-- Version: v11.9 SP6 11.9.6.7
-- File used only for Simulation

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Toplevel is

    port( AA            : in    std_logic;
          AB            : in    std_logic;
          ABSY          : in    std_logic;
          CLOCK         : in    std_logic;
          CU_SYNC       : in    std_logic;
          EMU_RX        : in    std_logic;
          FFU_EJECTED   : in    std_logic;
          FMC_CLK       : in    std_logic;
          FMC_NE1       : in    std_logic;
          FMC_NOE       : in    std_logic;
          RESET         : in    std_logic;
          TOP_UART_RX   : in    std_logic;
          UC_CONSOLE_EN : in    std_logic;
          UC_I2C4_SCL   : in    std_logic;
          UC_UART_TX    : in    std_logic;
          ACCE_SCL      : out   std_logic;
          ACLK          : out   std_logic;
          ACS           : out   std_logic;
          ACST          : out   std_logic;
          ARST          : out   std_logic;
          FMC_DA        : out   std_logic_vector(7 downto 0);
          FPGA_BUF_INT  : out   std_logic;
          FRAM_SCL      : out   std_logic;
          GYRO_SCL      : out   std_logic;
          L1WR          : out   std_logic;
          L2WR          : out   std_logic;
          L3WR          : out   std_logic;
          L4WR          : out   std_logic;
          LA0           : out   std_logic;
          LA1           : out   std_logic;
          LDCLK         : out   std_logic;
          LDCS          : out   std_logic;
          LDSDI         : out   std_logic;
          LED1          : out   std_logic;
          LED2          : out   std_logic;
          PRESSURE_SCL  : out   std_logic;
          SCIENCE_TX    : out   std_logic;
          TOP_UART_TX   : out   std_logic;
          UC_PWR_EN     : out   std_logic;
          UC_RESET      : out   std_logic;
          UC_UART_RX    : out   std_logic;
          ACCE_SDA      : inout std_logic := 'Z';
          FRAM_SDA      : inout std_logic := 'Z';
          GYRO_SDA      : inout std_logic := 'Z';
          PRESSURE_SDA  : inout std_logic := 'Z';
          UC_I2C4_SDA   : inout std_logic := 'Z'
        );

end Toplevel;

architecture DEF_ARCH of Toplevel is 

  component DFN1E1C1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN0E0C1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN0C1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AOI1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPAD_TRI
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN0P1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN0E1C1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOBI_IB_OB_EB
    port( D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          YIN  : in    std_logic := 'U';
          DOUT : out   std_logic;
          EOUT : out   std_logic;
          Y    : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPAD_BI
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic;
          PAD : inout   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOTRI_OB_EB
    port( D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          DOUT : out   std_logic;
          EOUT : out   std_logic
        );
  end component;

  component NAND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOIN_IB
    port( YIN : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM512X18
    generic (MEMORYFILE:string := "");

    port( RADDR8 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          WADDR8 : in    std_logic := 'U';
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          WD17   : in    std_logic := 'U';
          WD16   : in    std_logic := 'U';
          WD15   : in    std_logic := 'U';
          WD14   : in    std_logic := 'U';
          WD13   : in    std_logic := 'U';
          WD12   : in    std_logic := 'U';
          WD11   : in    std_logic := 'U';
          WD10   : in    std_logic := 'U';
          WD9    : in    std_logic := 'U';
          WD8    : in    std_logic := 'U';
          WD7    : in    std_logic := 'U';
          WD6    : in    std_logic := 'U';
          WD5    : in    std_logic := 'U';
          WD4    : in    std_logic := 'U';
          WD3    : in    std_logic := 'U';
          WD2    : in    std_logic := 'U';
          WD1    : in    std_logic := 'U';
          WD0    : in    std_logic := 'U';
          RW0    : in    std_logic := 'U';
          RW1    : in    std_logic := 'U';
          WW0    : in    std_logic := 'U';
          WW1    : in    std_logic := 'U';
          PIPE   : in    std_logic := 'U';
          REN    : in    std_logic := 'U';
          WEN    : in    std_logic := 'U';
          RCLK   : in    std_logic := 'U';
          WCLK   : in    std_logic := 'U';
          RESET  : in    std_logic := 'U';
          RD17   : out   std_logic;
          RD16   : out   std_logic;
          RD15   : out   std_logic;
          RD14   : out   std_logic;
          RD13   : out   std_logic;
          RD12   : out   std_logic;
          RD11   : out   std_logic;
          RD10   : out   std_logic;
          RD9    : out   std_logic;
          RD8    : out   std_logic;
          RD7    : out   std_logic;
          RD6    : out   std_logic;
          RD5    : out   std_logic;
          RD4    : out   std_logic;
          RD3    : out   std_logic;
          RD2    : out   std_logic;
          RD1    : out   std_logic;
          RD0    : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MIN3X
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0P1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFI1E1C1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          QN  : out   std_logic
        );
  end component;

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component AXO7
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MIN3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XAI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO16
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN0E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN0E0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AXO2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI7
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI4
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPAD_IN
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component AO18
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN0E0P1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXO5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ZOR3I
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1P1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AXO6
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port(Y : out std_logic); 
  end component;

  component VCC
    port(Y : out std_logic); 
  end component;

    signal CLKINT_0_Y_0, CLKINT_1_Y, CLKINT_2_Y, 
        ClockDivs_0_clk_800kHz, \SweepTable_0_RD[0]\, 
        \SweepTable_0_RD[1]\, \SweepTable_0_RD[2]\, 
        \SweepTable_0_RD[3]\, \SweepTable_0_RD[4]\, 
        \SweepTable_0_RD[5]\, \SweepTable_0_RD[6]\, 
        \SweepTable_0_RD[7]\, \SweepTable_0_RD[8]\, 
        \SweepTable_0_RD[9]\, \SweepTable_0_RD[10]\, 
        \SweepTable_0_RD[11]\, \SweepTable_0_RD[12]\, 
        \SweepTable_0_RD[13]\, \SweepTable_0_RD[14]\, 
        \SweepTable_0_RD[15]\, \SweepTable_1_RD[0]\, 
        \SweepTable_1_RD[1]\, \SweepTable_1_RD[2]\, 
        \SweepTable_1_RD[3]\, \SweepTable_1_RD[4]\, 
        \SweepTable_1_RD[5]\, \SweepTable_1_RD[6]\, 
        \SweepTable_1_RD[7]\, \SweepTable_1_RD[8]\, 
        \SweepTable_1_RD[9]\, \SweepTable_1_RD[10]\, 
        \SweepTable_1_RD[11]\, \SweepTable_1_RD[12]\, 
        \SweepTable_1_RD[13]\, \SweepTable_1_RD[14]\, 
        \SweepTable_1_RD[15]\, \General_Controller_0_st_wdata[0]\, 
        \General_Controller_0_st_wdata[1]\, 
        \General_Controller_0_st_wdata[2]\, 
        \General_Controller_0_st_wdata[3]\, 
        \General_Controller_0_st_wdata[4]\, 
        \General_Controller_0_st_wdata[5]\, 
        \General_Controller_0_st_wdata[6]\, 
        \General_Controller_0_st_wdata[7]\, 
        \General_Controller_0_st_wdata[8]\, 
        \General_Controller_0_st_wdata[9]\, 
        \General_Controller_0_st_wdata[10]\, 
        \General_Controller_0_st_wdata[11]\, 
        \General_Controller_0_st_wdata[12]\, 
        \General_Controller_0_st_wdata[13]\, 
        \General_Controller_0_st_wdata[14]\, 
        \General_Controller_0_st_wdata[15]\, 
        \General_Controller_0_st_waddr[0]\, 
        \General_Controller_0_st_waddr[1]\, 
        \General_Controller_0_st_waddr[2]\, 
        \General_Controller_0_st_waddr[3]\, 
        \General_Controller_0_st_waddr[4]\, 
        \General_Controller_0_st_waddr[5]\, 
        \General_Controller_0_st_waddr[6]\, 
        \General_Controller_0_st_waddr[7]\, 
        \TableSelect_0_RADDR[0]\, \TableSelect_0_RADDR[1]\, 
        \TableSelect_0_RADDR[2]\, \TableSelect_0_RADDR[3]\, 
        \TableSelect_0_RADDR[4]\, \TableSelect_0_RADDR[5]\, 
        \TableSelect_0_RADDR[6]\, \TableSelect_0_RADDR[7]\, 
        \SweepTable_1.WEBP\, \SweepTable_1.WEAP\, 
        \SweepTable_0.WEAP\, sda_cl_1_RNIGPAD, 
        \Sensors_0.Pressure_Sensor_0.I2C_Master_0.sda_1\, 
        sda_cl_1_RNITJT01, \Sensors_0.Gyro_0.I2C_Master_0.sda_1\, 
        sda_cl_1_RNIBFPP, 
        \Sensors_0.Accelerometer_0.I2C_Master_0.sda_1\, 
        \I2C_PassThrough_0.state[2]\, 
        \I2C_PassThrough_0.state[3]\, ACCE_SDA_in, FRAM_SDA_in, 
        GYRO_SDA_in, PRESSURE_SDA_in, UC_I2C4_SDA_in, AA_c, AB_c, 
        CLOCK_c, CU_SYNC_c, EMU_RX_c, FFU_EJECTED_c, FMC_CLK_c, 
        FMC_NOE_c, RESET_c, TOP_UART_RX_c, UC_CONSOLE_EN_c, 
        UC_UART_TX_c, ACCE_SCL_c, ACLK_c, ACS_c, ARST_c, 
        \FMC_DA_c[0]\, \FMC_DA_c[1]\, \FMC_DA_c[2]\, 
        \FMC_DA_c[3]\, \FMC_DA_c[4]\, \FMC_DA_c[5]\, 
        \FMC_DA_c[6]\, \FMC_DA_c[7]\, FPGA_BUF_INT_c, 
        FRAM_SCL_c_c, GYRO_SCL_c, L1WR_c, L2WR_c, L3WR_c, L4WR_c, 
        LA0_c, LA1_c, LDCLK_c, LDCS_c, LDSDI_c, LED1_c, LED2_c, 
        PRESSURE_SCL_c, SCIENCE_TX_c_c, UC_PWR_EN_c, UC_UART_RX_c, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[0]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[1]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[2]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[3]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[4]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[5]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[6]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[7]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[8]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[9]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[10]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[11]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[12]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[13]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[14]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[15]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[16]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[17]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[18]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[19]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[20]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[21]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[22]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[23]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[24]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[25]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[26]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[27]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[28]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[29]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[30]\, 
        \Data_Saving_0/Packet_Saver_0_data_out_0[31]\, 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[9]\, 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[0]\\\\\, 
        \VCC\, \GND\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[4]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[1]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[6]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[2]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[3]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[1]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[2]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[7]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[0]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[2]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[7]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/MEMWENEG\, 
        \Data_Saving_0/FPGA_Buffer_0/MEMRENEG\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[5]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[6]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[1]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[7]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[0]\\\\\, 
        \SweepTable_0/WEBP\, \GS_Readout_0/subState[0]_net_1\, 
        \GS_Readout_0/subState_0[0]\, \ClockDivs_0/clk_800kHz_i\, 
        \FMC_DA_pad[6]/U0/NET1\, \FMC_DA_pad[6]/U0/NET2\, 
        \LED1_pad/U0/NET1\, \LED1_pad/U0/NET2\, 
        \ACCE_SDA_pad/U0/NET1\, \ACCE_SDA_pad/U0/NET2\, 
        \ACCE_SDA_pad/U0/NET3\, \FMC_DA_pad[7]/U0/NET1\, 
        \FMC_DA_pad[7]/U0/NET2\, \UC_UART_TX_pad/U0/NET1\, 
        \UC_RESET_pad/U0/NET1\, \UC_RESET_pad/U0/NET2\, 
        \UC_PWR_EN_pad/U0/NET1\, \UC_PWR_EN_pad/U0/NET2\, 
        \FPGA_BUF_INT_pad/U0/NET1\, \FPGA_BUF_INT_pad/U0/NET2\, 
        \FRAM_SCL_pad/U0/NET1\, \FRAM_SCL_pad/U0/NET2\, 
        \CU_SYNC_pad/U0/NET1\, \CLOCK_pad/U0/NET1\, 
        \FMC_DA_pad[3]/U0/NET1\, \FMC_DA_pad[3]/U0/NET2\, 
        \ACCE_SCL_pad/U0/NET1\, \ACCE_SCL_pad/U0/NET2\, 
        \FMC_DA_pad[0]/U0/NET1\, \FMC_DA_pad[0]/U0/NET2\, 
        \RESET_pad/U0/NET1\, \LDCLK_pad/U0/NET1\, 
        \LDCLK_pad/U0/NET2\, \TOP_UART_TX_pad/U0/NET1\, 
        \TOP_UART_TX_pad/U0/NET2\, \UC_CONSOLE_EN_pad/U0/NET1\, 
        \FMC_DA_pad[1]/U0/NET1\, \FMC_DA_pad[1]/U0/NET2\, 
        \UC_I2C4_SCL_pad/U0/NET1\, \GYRO_SCL_pad/U0/NET1\, 
        \GYRO_SCL_pad/U0/NET2\, \TOP_UART_RX_pad/U0/NET1\, 
        \FMC_DA_pad[4]/U0/NET1\, \FMC_DA_pad[4]/U0/NET2\, 
        \ACLK_pad/U0/NET1\, \ACLK_pad/U0/NET2\, 
        \L4WR_pad/U0/NET1\, \L4WR_pad/U0/NET2\, 
        \LDSDI_pad/U0/NET1\, \LDSDI_pad/U0/NET2\, 
        \L1WR_pad/U0/NET1\, \L1WR_pad/U0/NET2\, \AA_pad/U0/NET1\, 
        \ACST_pad/U0/NET1\, \ACST_pad/U0/NET2\, 
        \EMU_RX_pad/U0/NET1\, \FMC_DA_pad[5]/U0/NET1\, 
        \FMC_DA_pad[5]/U0/NET2\, \LED2_pad/U0/NET1\, 
        \LED2_pad/U0/NET2\, \LA0_pad/U0/NET1\, \LA0_pad/U0/NET2\, 
        \AB_pad/U0/NET1\, \UC_UART_RX_pad/U0/NET1\, 
        \UC_UART_RX_pad/U0/NET2\, \L3WR_pad/U0/NET1\, 
        \L3WR_pad/U0/NET2\, \UC_I2C4_SDA_pad/U0/NET1\, 
        \UC_I2C4_SDA_pad/U0/NET2\, \UC_I2C4_SDA_pad/U0/NET3\, 
        \GYRO_SDA_pad/U0/NET1\, \GYRO_SDA_pad/U0/NET2\, 
        \GYRO_SDA_pad/U0/NET3\, \PRESSURE_SDA_pad/U0/NET1\, 
        \PRESSURE_SDA_pad/U0/NET2\, \PRESSURE_SDA_pad/U0/NET3\, 
        \FMC_CLK_pad/U0/NET1\, \FMC_NOE_pad/U0/NET1\, 
        \PRESSURE_SCL_pad/U0/NET1\, \PRESSURE_SCL_pad/U0/NET2\, 
        \SCIENCE_TX_pad/U0/NET1\, \SCIENCE_TX_pad/U0/NET2\, 
        \FFU_EJECTED_pad/U0/NET1\, \FMC_DA_pad[2]/U0/NET1\, 
        \FMC_DA_pad[2]/U0/NET2\, \LA1_pad/U0/NET1\, 
        \LA1_pad/U0/NET2\, \L2WR_pad/U0/NET1\, \L2WR_pad/U0/NET2\, 
        \LDCS_pad/U0/NET1\, \LDCS_pad/U0/NET2\, 
        \ARST_pad/U0/NET1\, \ARST_pad/U0/NET2\, 
        \FRAM_SDA_pad/U0/NET1\, \FRAM_SDA_pad/U0/NET2\, 
        \FRAM_SDA_pad/U0/NET3\, \ACS_pad/U0/NET1\, 
        \ACS_pad/U0/NET2\, \ClockDivs_0/cnt_800kHz[0]_net_1\, 
        \ClockDivs_0/cnt_800kHz[1]_net_1\, 
        \ClockDivs_0/cnt_800kHz[2]_net_1\, 
        \ClockDivs_0/cnt_800kHz[3]_net_1\, 
        \ClockDivs_0/cnt_800kHz[4]_net_1\, 
        \Communications_0/FFU_Command_Checker_0/state[0]_net_1\, 
        \Communications_0/FFU_Command_Checker_0/state[1]_net_1\, 
        \Communications_0/FFU_Command_Checker_0_rmu_oen\, 
        \Communications_0/UART_0/rx_byte[0]_net_1\, 
        \Communications_0/UART_0/rx_byte[1]_net_1\, 
        \Communications_0/UART_0/rx_byte[2]_net_1\, 
        \Communications_0/UART_0/rx_byte[3]_net_1\, 
        \Communications_0/UART_0/rx_byte[4]_net_1\, 
        \Communications_0/UART_0/rx_byte[5]_net_1\, 
        \Communications_0/UART_0/rx_byte[6]_net_1\, 
        \Communications_0/UART_0/rx_byte[7]_net_1\, 
        \Communications_0/UART_0/rx_clk_count[23]_net_1\, 
        \Communications_0/UART_0/rx_clk_count[24]_net_1\, 
        \Communications_0/UART_0/rx_clk_count[25]_net_1\, 
        \Communications_0/UART_0/rx_clk_count[26]_net_1\, 
        \Communications_0/UART_0/rx_clk_count[27]_net_1\, 
        \Communications_0/UART_0/rx_clk_count[28]_net_1\, 
        \Communications_0/UART_0/rx_clk_count[29]_net_1\, 
        \Communications_0/UART_0/rx_clk_count[30]_net_1\, 
        \Communications_0/UART_0/rx_clk_count_c0\, 
        \Communications_0/UART_0/rx_count[0]_net_1\, 
        \Communications_0/UART_0/rx_count[1]_net_1\, 
        \Communications_0/UART_0/rx_count[2]_net_1\, 
        \Communications_0/UART_0/rx_state[0]_net_1\, 
        \Communications_0/UART_0/rx_state[1]_net_1\, 
        \Communications_0/UART_0/tx_byte[0]_net_1\, 
        \Communications_0/UART_0/tx_byte[1]_net_1\, 
        \Communications_0/UART_0/tx_byte[2]_net_1\, 
        \Communications_0/UART_0/tx_byte[3]_net_1\, 
        \Communications_0/UART_0/tx_byte[4]_net_1\, 
        \Communications_0/UART_0/tx_byte[5]_net_1\, 
        \Communications_0/UART_0/tx_byte[6]_net_1\, 
        \Communications_0/UART_0/tx_byte[7]_net_1\, 
        \Communications_0/UART_0/tx_clk_count[0]_net_1\, 
        \Communications_0/UART_0/tx_clk_count[1]_net_1\, 
        \Communications_0/UART_0/tx_clk_count_i_0[2]\, 
        \Communications_0/UART_0/tx_clk_count_i_0[3]\, 
        \Communications_0/UART_0/tx_clk_count_i_0[4]\, 
        \Communications_0/UART_0/tx_clk_count_i_0[5]\, 
        \Communications_0/UART_0/tx_clk_count_i_0[6]\, 
        \Communications_0/UART_0/tx_clk_count_i_0[7]\, 
        \Communications_0/UART_0/tx_clk_count_i_0[8]\, 
        \Communications_0/UART_0/tx_count[0]_net_1\, 
        \Communications_0/UART_0/tx_count[1]_net_1\, 
        \Communications_0/UART_0/tx_count[2]_net_1\, 
        \Communications_0/UART_0/tx_state[0]_net_1\, 
        \Communications_0/UART_0/tx_state[1]_net_1\, 
        \Communications_0/UART_0_recv[0]\, 
        \Communications_0/UART_0_recv[1]\, 
        \Communications_0/UART_0_recv[2]\, 
        \Communications_0/UART_0_recv[3]\, 
        \Communications_0/UART_0_recv[4]\, 
        \Communications_0/UART_0_recv[5]\, 
        \Communications_0/UART_0_recv[6]\, 
        \Communications_0/UART_0_recv[7]\, 
        \Communications_0/UART_0_rx_rdy\, 
        \Communications_0/UART_0_tx\, 
        \Communications_0/UART_1/rx_byte[0]_net_1\, 
        \Communications_0/UART_1/rx_byte[1]_net_1\, 
        \Communications_0/UART_1/rx_byte[2]_net_1\, 
        \Communications_0/UART_1/rx_byte[3]_net_1\, 
        \Communications_0/UART_1/rx_byte[4]_net_1\, 
        \Communications_0/UART_1/rx_byte[5]_net_1\, 
        \Communications_0/UART_1/rx_byte[6]_net_1\, 
        \Communications_0/UART_1/rx_byte[7]_net_1\, 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\, 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\, 
        \Communications_0/UART_1/rx_clk_count[25]_net_1\, 
        \Communications_0/UART_1/rx_clk_count[26]_net_1\, 
        \Communications_0/UART_1/rx_clk_count[27]_net_1\, 
        \Communications_0/UART_1/rx_clk_count[28]_net_1\, 
        \Communications_0/UART_1/rx_clk_count[29]_net_1\, 
        \Communications_0/UART_1/rx_clk_count[30]_net_1\, 
        \Communications_0/UART_1/rx_clk_count_c0\, 
        \Communications_0/UART_1/rx_count[0]_net_1\, 
        \Communications_0/UART_1/rx_count[1]_net_1\, 
        \Communications_0/UART_1/rx_count[2]_net_1\, 
        \Communications_0/UART_1/rx_state[0]_net_1\, 
        \Communications_0/UART_1/rx_state[1]_net_1\, 
        \Communications_0/UART_1/tx_byte[0]_net_1\, 
        \Communications_0/UART_1/tx_byte[1]_net_1\, 
        \Communications_0/UART_1/tx_byte[2]_net_1\, 
        \Communications_0/UART_1/tx_byte[3]_net_1\, 
        \Communications_0/UART_1/tx_byte[4]_net_1\, 
        \Communications_0/UART_1/tx_byte[5]_net_1\, 
        \Communications_0/UART_1/tx_byte[6]_net_1\, 
        \Communications_0/UART_1/tx_byte[7]_net_1\, 
        \Communications_0/UART_1/tx_clk_count[0]_net_1\, 
        \Communications_0/UART_1/tx_clk_count[1]_net_1\, 
        \Communications_0/UART_1/tx_clk_count_i_0[2]\, 
        \Communications_0/UART_1/tx_clk_count_i_0[3]\, 
        \Communications_0/UART_1/tx_clk_count_i_0[4]\, 
        \Communications_0/UART_1/tx_clk_count_i_0[5]\, 
        \Communications_0/UART_1/tx_clk_count_i_0[6]\, 
        \Communications_0/UART_1/tx_clk_count_i_0[7]\, 
        \Communications_0/UART_1/tx_clk_count_i_0[8]\, 
        \Communications_0/UART_1/tx_count[0]_net_1\, 
        \Communications_0/UART_1/tx_count[1]_net_1\, 
        \Communications_0/UART_1/tx_count[2]_net_1\, 
        \Communications_0/UART_1/tx_state[0]_net_1\, 
        \Communications_0/UART_1/tx_state[1]_net_1\, 
        \Communications_0/UART_1_tx\, 
        \Communications_0_ext_recv[0]\, 
        \Communications_0_ext_recv[1]\, 
        \Communications_0_ext_recv[2]\, 
        \Communications_0_ext_recv[3]\, 
        \Communications_0_ext_recv[4]\, 
        \Communications_0_ext_recv[5]\, 
        \Communications_0_ext_recv[6]\, 
        \Communications_0_ext_recv[7]\, 
        Communications_0_ext_rx_rdy, Communications_0_ext_tx_rdy, 
        \Communications_0_uc_recv[0]\, 
        \Communications_0_uc_recv[1]\, 
        \Communications_0_uc_recv[2]\, 
        \Communications_0_uc_recv[3]\, 
        \Communications_0_uc_recv[4]\, 
        \Communications_0_uc_recv[5]\, 
        \Communications_0_uc_recv[6]\, 
        \Communications_0_uc_recv[7]\, Communications_0_uc_rx_rdy, 
        Communications_0_uc_tx_rdy, 
        \Data_Hub_Packets_0_status_packet[0]\, 
        \Data_Hub_Packets_0_status_packet[1]\, 
        \Data_Hub_Packets_0_status_packet[2]\, 
        \Data_Hub_Packets_0_status_packet[3]\, 
        \Data_Hub_Packets_0_status_packet[40]\, 
        \Data_Hub_Packets_0_status_packet[41]\, 
        \Data_Hub_Packets_0_status_packet[42]\, 
        \Data_Hub_Packets_0_status_packet[43]\, 
        \Data_Hub_Packets_0_status_packet[44]\, 
        \Data_Hub_Packets_0_status_packet[45]\, 
        \Data_Hub_Packets_0_status_packet[46]\, 
        \Data_Hub_Packets_0_status_packet[47]\, 
        \Data_Hub_Packets_0_status_packet[48]\, 
        \Data_Hub_Packets_0_status_packet[49]\, 
        \Data_Hub_Packets_0_status_packet[4]\, 
        \Data_Hub_Packets_0_status_packet[50]\, 
        \Data_Hub_Packets_0_status_packet[51]\, 
        \Data_Hub_Packets_0_status_packet[52]\, 
        \Data_Hub_Packets_0_status_packet[53]\, 
        \Data_Hub_Packets_0_status_packet[54]\, 
        \Data_Hub_Packets_0_status_packet[55]\, 
        \Data_Hub_Packets_0_status_packet[56]\, 
        \Data_Hub_Packets_0_status_packet[57]\, 
        \Data_Hub_Packets_0_status_packet[58]\, 
        \Data_Hub_Packets_0_status_packet[59]\, 
        \Data_Hub_Packets_0_status_packet[5]\, 
        \Data_Hub_Packets_0_status_packet[60]\, 
        \Data_Hub_Packets_0_status_packet[61]\, 
        \Data_Hub_Packets_0_status_packet[62]\, 
        \Data_Hub_Packets_0_status_packet[63]\, 
        \Data_Hub_Packets_0_status_packet[6]\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_10_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_11_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_12_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_13_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_14_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_15_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_16_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_17_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_18_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_19_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_1_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_20_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_2_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_3_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_4_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_5_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_6_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_7_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_8_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_9_Q\, 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\, 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[10]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[8]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[10]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[2]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[3]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[4]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[5]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[6]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[7]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[8]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[9]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[10]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[2]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[3]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[4]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[5]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[6]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[7]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[8]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[9]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[0]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[1]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[2]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[3]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[4]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[5]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[6]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[7]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[8]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[0]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[1]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[2]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[3]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[4]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[5]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[6]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[7]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[8]\\\\\, 
        \Data_Saving_0/FPGA_Buffer_0/empty\, 
        \Data_Saving_0/FPGA_Buffer_0/full\, 
        \Data_Saving_0/FPGA_Buffer_0_afull\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[0]_net_1\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[1]_net_1\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[2]_net_1\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[3]_net_1\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[4]_net_1\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[5]_net_1\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[6]_net_1\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[7]_net_1\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[8]_net_1\, 
        \Data_Saving_0/Interrupt_Generator_0/counter[9]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/acc_flag_net_1\, 
        \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\, 
        \Data_Saving_0/Packet_Saver_0/gyro_flag_net_1\, 
        \Data_Saving_0/Packet_Saver_0/mag_flag_net_1\, 
        \Data_Saving_0/Packet_Saver_0/old_acc_new_data_i_0\, 
        \Data_Saving_0/Packet_Saver_0/old_ch_0_new_data_i_0\, 
        \Data_Saving_0/Packet_Saver_0/old_gyro_new_data_i_0\, 
        \Data_Saving_0/Packet_Saver_0/old_mag_new_data_i_0\, 
        \Data_Saving_0/Packet_Saver_0/old_pressure_new_data_i_0\, 
        \Data_Saving_0/Packet_Saver_0/old_status_new_data_i_0\, 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/pressure_flag_net_1\, 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/status_flag_net_1\, 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/word_cnt[1]_net_1\, 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, 
        \Data_Saving_0/Packet_Saver_0_we\, 
        \Eject_Signal_Debounce_0/ms_cnt[0]_net_1\, 
        \Eject_Signal_Debounce_0/ms_cnt[1]_net_1\, 
        \Eject_Signal_Debounce_0/ms_cnt[2]_net_1\, 
        \Eject_Signal_Debounce_0/ms_cnt[3]_net_1\, 
        \Eject_Signal_Debounce_0/ms_cnt[4]_net_1\, 
        \Eject_Signal_Debounce_0/ms_cnt[5]_net_1\, 
        \Eject_Signal_Debounce_0/old_1kHz_i_0\, 
        \Eject_Signal_Debounce_0/state[0]_net_1\, 
        \Eject_Signal_Debounce_0/state[1]_net_1\, 
        Eject_Signal_Debounce_0_ffu_ejected_out, 
        \GS_Readout_0/prevState[0]_net_1\, 
        \GS_Readout_0/prevState[1]_net_1\, 
        \GS_Readout_0/prevState[2]_net_1\, 
        \GS_Readout_0/prevState[3]_net_1\, 
        \GS_Readout_0/prevState[4]_net_1\, 
        \GS_Readout_0/prevState[5]_net_1\, 
        \GS_Readout_0/prevState[7]_net_1\, 
        \GS_Readout_0/state[0]_net_1\, 
        \GS_Readout_0/state[1]_net_1\, 
        \GS_Readout_0/state[2]_net_1\, 
        \GS_Readout_0/state[3]_net_1\, 
        \GS_Readout_0/state[4]_net_1\, 
        \GS_Readout_0/state[5]_net_1\, 
        \GS_Readout_0/state[6]_net_1\, 
        \GS_Readout_0/state[7]_net_1\, 
        \GS_Readout_0/subState[1]_net_1\, 
        \GS_Readout_0/subState[2]_net_1\, 
        \GS_Readout_0/subState[3]_net_1\, 
        \GS_Readout_0/subState[4]_net_1\, \GS_Readout_0_send[0]\, 
        \GS_Readout_0_send[1]\, \GS_Readout_0_send[2]\, 
        \GS_Readout_0_send[3]\, \GS_Readout_0_send[4]\, 
        \GS_Readout_0_send[5]\, \GS_Readout_0_send[6]\, 
        \GS_Readout_0_send[7]\, GS_Readout_0_wen, 
        \General_Controller_0/command[0]_net_1\, 
        \General_Controller_0/command[1]_net_1\, 
        \General_Controller_0/command[2]_net_1\, 
        \General_Controller_0/command[3]_net_1\, 
        \General_Controller_0/command[4]_net_1\, 
        \General_Controller_0/command[5]_net_1\, 
        \General_Controller_0/command[6]_net_1\, 
        \General_Controller_0/command[7]_net_1\, 
        \General_Controller_0/constant_bias_probe_id[0]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[0]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[10]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[11]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[12]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[13]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[14]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[15]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[1]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[2]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[3]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[4]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[5]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[6]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[7]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[8]_net_1\, 
        \General_Controller_0/constant_bias_voltage_0[9]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[0]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[10]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[11]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[12]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[13]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[14]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[15]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[1]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[2]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[3]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[4]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[5]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[6]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[7]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[8]_net_1\, 
        \General_Controller_0/constant_bias_voltage_1[9]_net_1\, 
        \General_Controller_0/ext_rx_state[0]_net_1\, 
        \General_Controller_0/ext_rx_state_i_0[1]\, 
        \General_Controller_0/flight_state[0]_net_1\, 
        \General_Controller_0/flight_state[1]_net_1\, 
        \General_Controller_0/flight_state[2]_net_1\, 
        \General_Controller_0/flight_state[3]_net_1\, 
        \General_Controller_0/flight_state[4]_net_1\, 
        \General_Controller_0/mission_mode_net_1\, 
        \General_Controller_0/old_1Hz_i_0\, 
        \General_Controller_0/old_status_packet_clk_i_0\, 
        \General_Controller_0/state_seconds[0]_net_1\, 
        \General_Controller_0/state_seconds[10]_net_1\, 
        \General_Controller_0/state_seconds[11]_net_1\, 
        \General_Controller_0/state_seconds[12]_net_1\, 
        \General_Controller_0/state_seconds[13]_net_1\, 
        \General_Controller_0/state_seconds[14]_net_1\, 
        \General_Controller_0/state_seconds[15]_net_1\, 
        \General_Controller_0/state_seconds[16]_net_1\, 
        \General_Controller_0/state_seconds[17]_net_1\, 
        \General_Controller_0/state_seconds[18]_net_1\, 
        \General_Controller_0/state_seconds[19]_net_1\, 
        \General_Controller_0/state_seconds[1]_net_1\, 
        \General_Controller_0/state_seconds[2]_net_1\, 
        \General_Controller_0/state_seconds[3]_net_1\, 
        \General_Controller_0/state_seconds[4]_net_1\, 
        \General_Controller_0/state_seconds[5]_net_1\, 
        \General_Controller_0/state_seconds[6]_net_1\, 
        \General_Controller_0/state_seconds[7]_net_1\, 
        \General_Controller_0/state_seconds[8]_net_1\, 
        \General_Controller_0/state_seconds[9]_net_1\, 
        \General_Controller_0/sweep_table_nof_steps[0]_net_1\, 
        \General_Controller_0/sweep_table_nof_steps[1]_net_1\, 
        \General_Controller_0/sweep_table_nof_steps[2]_net_1\, 
        \General_Controller_0/sweep_table_nof_steps[3]_net_1\, 
        \General_Controller_0/sweep_table_nof_steps[4]_net_1\, 
        \General_Controller_0/sweep_table_nof_steps[5]_net_1\, 
        \General_Controller_0/sweep_table_nof_steps[6]_net_1\, 
        \General_Controller_0/sweep_table_nof_steps[7]_net_1\, 
        \General_Controller_0/sweep_table_points[0]_net_1\, 
        \General_Controller_0/sweep_table_points[10]_net_1\, 
        \General_Controller_0/sweep_table_points[11]_net_1\, 
        \General_Controller_0/sweep_table_points[12]_net_1\, 
        \General_Controller_0/sweep_table_points[13]_net_1\, 
        \General_Controller_0/sweep_table_points[14]_net_1\, 
        \General_Controller_0/sweep_table_points[15]_net_1\, 
        \General_Controller_0/sweep_table_points[1]_net_1\, 
        \General_Controller_0/sweep_table_points[2]_net_1\, 
        \General_Controller_0/sweep_table_points[3]_net_1\, 
        \General_Controller_0/sweep_table_points[4]_net_1\, 
        \General_Controller_0/sweep_table_points[5]_net_1\, 
        \General_Controller_0/sweep_table_points[6]_net_1\, 
        \General_Controller_0/sweep_table_points[7]_net_1\, 
        \General_Controller_0/sweep_table_points[8]_net_1\, 
        \General_Controller_0/sweep_table_points[9]_net_1\, 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, 
        \General_Controller_0/sweep_table_probe_id[1]_net_1\, 
        \General_Controller_0/sweep_table_probe_id[2]_net_1\, 
        \General_Controller_0/sweep_table_probe_id[3]_net_1\, 
        \General_Controller_0/sweep_table_probe_id[4]_net_1\, 
        \General_Controller_0/sweep_table_probe_id[5]_net_1\, 
        \General_Controller_0/sweep_table_probe_id[6]_net_1\, 
        \General_Controller_0/sweep_table_probe_id[7]_net_1\, 
        \General_Controller_0/sweep_table_read_value[0]_net_1\, 
        \General_Controller_0/sweep_table_read_value[10]_net_1\, 
        \General_Controller_0/sweep_table_read_value[11]_net_1\, 
        \General_Controller_0/sweep_table_read_value[12]_net_1\, 
        \General_Controller_0/sweep_table_read_value[13]_net_1\, 
        \General_Controller_0/sweep_table_read_value[14]_net_1\, 
        \General_Controller_0/sweep_table_read_value[15]_net_1\, 
        \General_Controller_0/sweep_table_read_value[1]_net_1\, 
        \General_Controller_0/sweep_table_read_value[2]_net_1\, 
        \General_Controller_0/sweep_table_read_value[3]_net_1\, 
        \General_Controller_0/sweep_table_read_value[4]_net_1\, 
        \General_Controller_0/sweep_table_read_value[5]_net_1\, 
        \General_Controller_0/sweep_table_read_value[6]_net_1\, 
        \General_Controller_0/sweep_table_read_value[7]_net_1\, 
        \General_Controller_0/sweep_table_read_value[8]_net_1\, 
        \General_Controller_0/sweep_table_read_value[9]_net_1\, 
        \General_Controller_0/sweep_table_read_wait[30]_net_1\, 
        \General_Controller_0/sweep_table_read_wait[31]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[0]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[10]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[11]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[12]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[13]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[14]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[15]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[1]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[2]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[3]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[4]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[5]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[6]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[7]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[8]_net_1\, 
        \General_Controller_0/sweep_table_sample_skip[9]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[0]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[10]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[11]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[12]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[13]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[14]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[15]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[1]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[2]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[3]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[4]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[5]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[6]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[7]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[8]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_point[9]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[0]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[10]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[11]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[12]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[13]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[14]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[15]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[1]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[2]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[3]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[4]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[5]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[6]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[7]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[8]_net_1\, 
        \General_Controller_0/sweep_table_samples_per_step[9]_net_1\, 
        \General_Controller_0/sweep_table_step_id[0]_net_1\, 
        \General_Controller_0/sweep_table_step_id[1]_net_1\, 
        \General_Controller_0/sweep_table_step_id[2]_net_1\, 
        \General_Controller_0/sweep_table_step_id[3]_net_1\, 
        \General_Controller_0/sweep_table_step_id[4]_net_1\, 
        \General_Controller_0/sweep_table_step_id[5]_net_1\, 
        \General_Controller_0/sweep_table_step_id[6]_net_1\, 
        \General_Controller_0/sweep_table_step_id[7]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[0]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[10]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[11]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[12]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[13]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[14]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[15]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[1]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[2]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[3]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[4]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[5]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[6]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[7]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[8]_net_1\, 
        \General_Controller_0/sweep_table_sweep_cnt[9]_net_1\, 
        \General_Controller_0/sweep_table_write_value[0]_net_1\, 
        \General_Controller_0/sweep_table_write_value[10]_net_1\, 
        \General_Controller_0/sweep_table_write_value[11]_net_1\, 
        \General_Controller_0/sweep_table_write_value[12]_net_1\, 
        \General_Controller_0/sweep_table_write_value[13]_net_1\, 
        \General_Controller_0/sweep_table_write_value[14]_net_1\, 
        \General_Controller_0/sweep_table_write_value[15]_net_1\, 
        \General_Controller_0/sweep_table_write_value[1]_net_1\, 
        \General_Controller_0/sweep_table_write_value[2]_net_1\, 
        \General_Controller_0/sweep_table_write_value[3]_net_1\, 
        \General_Controller_0/sweep_table_write_value[4]_net_1\, 
        \General_Controller_0/sweep_table_write_value[5]_net_1\, 
        \General_Controller_0/sweep_table_write_value[6]_net_1\, 
        \General_Controller_0/sweep_table_write_value[7]_net_1\, 
        \General_Controller_0/sweep_table_write_value[8]_net_1\, 
        \General_Controller_0/sweep_table_write_value[9]_net_1\, 
        \General_Controller_0/sweep_table_write_wait[0]_net_1\, 
        \General_Controller_0/sweep_table_write_wait[1]_net_1\, 
        \General_Controller_0/temp_first_byte[0]_net_1\, 
        \General_Controller_0/temp_first_byte[1]_net_1\, 
        \General_Controller_0/temp_first_byte[2]_net_1\, 
        \General_Controller_0/temp_first_byte[3]_net_1\, 
        \General_Controller_0/temp_first_byte[4]_net_1\, 
        \General_Controller_0/temp_first_byte[5]_net_1\, 
        \General_Controller_0/temp_first_byte[6]_net_1\, 
        \General_Controller_0/temp_first_byte[7]_net_1\, 
        \General_Controller_0/uc_rx_byte[0]_net_1\, 
        \General_Controller_0/uc_rx_byte[1]_net_1\, 
        \General_Controller_0/uc_rx_byte[2]_net_1\, 
        \General_Controller_0/uc_rx_byte[3]_net_1\, 
        \General_Controller_0/uc_rx_byte[4]_net_1\, 
        \General_Controller_0/uc_rx_byte[5]_net_1\, 
        \General_Controller_0/uc_rx_byte[6]_net_1\, 
        \General_Controller_0/uc_rx_byte[7]_net_1\, 
        \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        \General_Controller_0/uc_rx_prev_state[0]_net_1\, 
        \General_Controller_0/uc_rx_prev_state[1]_net_1\, 
        \General_Controller_0/uc_rx_prev_state[2]_net_1\, 
        \General_Controller_0/uc_rx_prev_state[3]_net_1\, 
        \General_Controller_0/uc_rx_prev_state[4]_net_1\, 
        \General_Controller_0/uc_rx_state[0]_net_1\, 
        \General_Controller_0/uc_rx_state[1]_net_1\, 
        \General_Controller_0/uc_rx_state[2]_net_1\, 
        \General_Controller_0/uc_rx_state[3]_net_1\, 
        \General_Controller_0/uc_rx_state[4]_net_1\, 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        \General_Controller_0/uc_rx_state_0[1]_net_1\, 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, 
        \General_Controller_0/uc_rx_substate[0]_net_1\, 
        \General_Controller_0/uc_rx_substate[1]_net_1\, 
        \General_Controller_0/uc_rx_substate[2]_net_1\, 
        \General_Controller_0/uc_rx_substate[3]_net_1\, 
        \General_Controller_0/uc_rx_substate[4]_net_1\, 
        \General_Controller_0/uc_tx_nextstate[0]_net_1\, 
        \General_Controller_0/uc_tx_nextstate[1]_net_1\, 
        \General_Controller_0/uc_tx_nextstate[2]_net_1\, 
        \General_Controller_0/uc_tx_nextstate[3]_net_1\, 
        \General_Controller_0/uc_tx_nextstate[4]_net_1\, 
        \General_Controller_0/uc_tx_nextstate[5]_net_1\, 
        \General_Controller_0/uc_tx_nextstate[6]_net_1\, 
        \General_Controller_0/uc_tx_nextstate[7]_net_1\, 
        \General_Controller_0/uc_tx_state[0]_net_1\, 
        \General_Controller_0/uc_tx_state[12]_net_1\, 
        \General_Controller_0/uc_tx_state[14]_net_1\, 
        \General_Controller_0/uc_tx_state[15]_net_1\, 
        \General_Controller_0/uc_tx_state[1]_net_1\, 
        \General_Controller_0/uc_tx_state[2]_net_1\, 
        \General_Controller_0/uc_tx_state[3]_net_1\, 
        \General_Controller_0/uc_tx_state[4]_net_1\, 
        \General_Controller_0/uc_tx_state[5]_net_1\, 
        \General_Controller_0/uc_tx_state[6]_net_1\, 
        \General_Controller_0/uc_tx_state[7]_net_1\, 
        \General_Controller_0/uc_tx_substate[0]_net_1\, 
        \General_Controller_0/uc_tx_substate[1]_net_1\, 
        \General_Controller_0/uc_tx_substate[2]_net_1\, 
        \General_Controller_0/uc_tx_substate[3]_net_1\, 
        \General_Controller_0/uc_tx_substate[4]_net_1\, 
        \General_Controller_0/un10_uc_tx_rdy_i[1]\, 
        \General_Controller_0/un10_uc_tx_rdy_i[2]\, 
        \General_Controller_0/un10_uc_tx_rdy_i[3]\, 
        \General_Controller_0/un10_uc_tx_rdy_i[4]\, 
        \General_Controller_0/un10_uc_tx_rdy_i[5]\, 
        \General_Controller_0/un10_uc_tx_rdy_i[6]\, 
        \General_Controller_0/un10_uc_tx_rdy_i[7]\, 
        General_Controller_0_en_data_saving, 
        General_Controller_0_en_science_packets, 
        General_Controller_0_en_sensors, 
        General_Controller_0_exp_adc_reset, 
        General_Controller_0_ext_oen, 
        \General_Controller_0_gs_id[0]\, 
        \General_Controller_0_gs_id[1]\, 
        \General_Controller_0_gs_id[2]\, 
        \General_Controller_0_gs_id[3]\, 
        \General_Controller_0_gs_id[4]\, 
        \General_Controller_0_gs_id[5]\, 
        \General_Controller_0_gs_id[6]\, 
        \General_Controller_0_gs_id[7]\, 
        General_Controller_0_readout_en, 
        \General_Controller_0_st_raddr_1[0]\, 
        \General_Controller_0_st_raddr_1[1]\, 
        \General_Controller_0_st_raddr_1[2]\, 
        \General_Controller_0_st_raddr_1[3]\, 
        \General_Controller_0_st_raddr_1[4]\, 
        \General_Controller_0_st_raddr_1[5]\, 
        \General_Controller_0_st_raddr_1[6]\, 
        \General_Controller_0_st_raddr_1[7]\, 
        General_Controller_0_st_ren1, 
        General_Controller_0_status_new_data, 
        General_Controller_0_uc_oen, 
        \General_Controller_0_uc_send[0]\, 
        \General_Controller_0_uc_send[1]\, 
        \General_Controller_0_uc_send[2]\, 
        \General_Controller_0_uc_send[3]\, 
        \General_Controller_0_uc_send[4]\, 
        \General_Controller_0_uc_send[5]\, 
        \General_Controller_0_uc_send[6]\, 
        \General_Controller_0_uc_send[7]\, 
        General_Controller_0_uc_wen, 
        \General_Controller_0_unit_id[0]\, 
        \General_Controller_0_unit_id[1]\, 
        \General_Controller_0_unit_id[2]\, 
        \General_Controller_0_unit_id[3]\, 
        \General_Controller_0_unit_id[4]\, 
        \General_Controller_0_unit_id[5]\, 
        \General_Controller_0_unit_id[6]\, 
        \General_Controller_0_unit_id[7]\, HIEFFPLA_NET_0_71968, 
        HIEFFPLA_NET_0_71969, HIEFFPLA_NET_0_71970, 
        HIEFFPLA_NET_0_71971, HIEFFPLA_NET_0_71972, 
        HIEFFPLA_NET_0_71973, HIEFFPLA_NET_0_71974, 
        HIEFFPLA_NET_0_71975, HIEFFPLA_NET_0_71976, 
        HIEFFPLA_NET_0_71977, HIEFFPLA_NET_0_71978, 
        HIEFFPLA_NET_0_71979, HIEFFPLA_NET_0_71980, 
        HIEFFPLA_NET_0_71981, HIEFFPLA_NET_0_71982, 
        HIEFFPLA_NET_0_71983, HIEFFPLA_NET_0_71984, 
        HIEFFPLA_NET_0_71985, HIEFFPLA_NET_0_71986, 
        HIEFFPLA_NET_0_71987, HIEFFPLA_NET_0_71988, 
        HIEFFPLA_NET_0_71989, HIEFFPLA_NET_0_71990, 
        HIEFFPLA_NET_0_71991, HIEFFPLA_NET_0_71992, 
        HIEFFPLA_NET_0_71993, HIEFFPLA_NET_0_71994, 
        HIEFFPLA_NET_0_71995, HIEFFPLA_NET_0_71996, 
        HIEFFPLA_NET_0_71997, HIEFFPLA_NET_0_71998, 
        HIEFFPLA_NET_0_71999, HIEFFPLA_NET_0_72000, 
        HIEFFPLA_NET_0_72001, HIEFFPLA_NET_0_72002, 
        HIEFFPLA_NET_0_72003, HIEFFPLA_NET_0_72004, 
        HIEFFPLA_NET_0_72005, HIEFFPLA_NET_0_72006, 
        HIEFFPLA_NET_0_72007, HIEFFPLA_NET_0_72008, 
        HIEFFPLA_NET_0_72009, HIEFFPLA_NET_0_72010, 
        HIEFFPLA_NET_0_72011, HIEFFPLA_NET_0_72012, 
        HIEFFPLA_NET_0_72013, HIEFFPLA_NET_0_72014, 
        HIEFFPLA_NET_0_72015, HIEFFPLA_NET_0_72016, 
        HIEFFPLA_NET_0_72017, HIEFFPLA_NET_0_72018, 
        HIEFFPLA_NET_0_72019, HIEFFPLA_NET_0_72020, 
        HIEFFPLA_NET_0_72021, HIEFFPLA_NET_0_72022, 
        HIEFFPLA_NET_0_72023, HIEFFPLA_NET_0_72024, 
        HIEFFPLA_NET_0_72025, HIEFFPLA_NET_0_72026, 
        HIEFFPLA_NET_0_72027, HIEFFPLA_NET_0_72028, 
        HIEFFPLA_NET_0_72029, HIEFFPLA_NET_0_72030, 
        HIEFFPLA_NET_0_72031, HIEFFPLA_NET_0_72032, 
        HIEFFPLA_NET_0_72033, HIEFFPLA_NET_0_72034, 
        HIEFFPLA_NET_0_72035, HIEFFPLA_NET_0_72036, 
        HIEFFPLA_NET_0_72037, HIEFFPLA_NET_0_72038, 
        HIEFFPLA_NET_0_72039, HIEFFPLA_NET_0_72040, 
        HIEFFPLA_NET_0_72041, HIEFFPLA_NET_0_72042, 
        HIEFFPLA_NET_0_72043, HIEFFPLA_NET_0_72044, 
        HIEFFPLA_NET_0_72045, HIEFFPLA_NET_0_72046, 
        HIEFFPLA_NET_0_72047, HIEFFPLA_NET_0_72048, 
        HIEFFPLA_NET_0_72049, HIEFFPLA_NET_0_72050, 
        HIEFFPLA_NET_0_72051, HIEFFPLA_NET_0_72052, 
        HIEFFPLA_NET_0_72053, HIEFFPLA_NET_0_72054, 
        HIEFFPLA_NET_0_72055, HIEFFPLA_NET_0_72056, 
        HIEFFPLA_NET_0_72057, HIEFFPLA_NET_0_72058, 
        HIEFFPLA_NET_0_72059, HIEFFPLA_NET_0_72060, 
        HIEFFPLA_NET_0_72061, HIEFFPLA_NET_0_72062, 
        HIEFFPLA_NET_0_72063, HIEFFPLA_NET_0_72064, 
        HIEFFPLA_NET_0_72065, HIEFFPLA_NET_0_72066, 
        HIEFFPLA_NET_0_72067, HIEFFPLA_NET_0_72068, 
        HIEFFPLA_NET_0_72069, HIEFFPLA_NET_0_72070, 
        HIEFFPLA_NET_0_72071, HIEFFPLA_NET_0_72072, 
        HIEFFPLA_NET_0_72073, HIEFFPLA_NET_0_72074, 
        HIEFFPLA_NET_0_72075, HIEFFPLA_NET_0_72076, 
        HIEFFPLA_NET_0_72077, HIEFFPLA_NET_0_72078, 
        HIEFFPLA_NET_0_72079, HIEFFPLA_NET_0_72080, 
        HIEFFPLA_NET_0_72081, HIEFFPLA_NET_0_72082, 
        HIEFFPLA_NET_0_72083, HIEFFPLA_NET_0_72084, 
        HIEFFPLA_NET_0_72085, HIEFFPLA_NET_0_72086, 
        HIEFFPLA_NET_0_72087, HIEFFPLA_NET_0_72088, 
        HIEFFPLA_NET_0_72089, HIEFFPLA_NET_0_72090, 
        HIEFFPLA_NET_0_72091, HIEFFPLA_NET_0_72092, 
        HIEFFPLA_NET_0_72093, HIEFFPLA_NET_0_72094, 
        HIEFFPLA_NET_0_72095, HIEFFPLA_NET_0_72096, 
        HIEFFPLA_NET_0_72097, HIEFFPLA_NET_0_72098, 
        HIEFFPLA_NET_0_72099, HIEFFPLA_NET_0_72100, 
        HIEFFPLA_NET_0_72101, HIEFFPLA_NET_0_72102, 
        HIEFFPLA_NET_0_72103, HIEFFPLA_NET_0_72104, 
        HIEFFPLA_NET_0_72105, HIEFFPLA_NET_0_72106, 
        HIEFFPLA_NET_0_72107, HIEFFPLA_NET_0_72108, 
        HIEFFPLA_NET_0_72109, HIEFFPLA_NET_0_72110, 
        HIEFFPLA_NET_0_72111, HIEFFPLA_NET_0_72112, 
        HIEFFPLA_NET_0_72113, HIEFFPLA_NET_0_72114, 
        HIEFFPLA_NET_0_72115, HIEFFPLA_NET_0_72116, 
        HIEFFPLA_NET_0_72117, HIEFFPLA_NET_0_72118, 
        HIEFFPLA_NET_0_72119, HIEFFPLA_NET_0_72120, 
        HIEFFPLA_NET_0_72121, HIEFFPLA_NET_0_72122, 
        HIEFFPLA_NET_0_72123, HIEFFPLA_NET_0_72124, 
        HIEFFPLA_NET_0_72125, HIEFFPLA_NET_0_72126, 
        HIEFFPLA_NET_0_72127, HIEFFPLA_NET_0_72128, 
        HIEFFPLA_NET_0_72129, HIEFFPLA_NET_0_72130, 
        HIEFFPLA_NET_0_72131, HIEFFPLA_NET_0_72132, 
        HIEFFPLA_NET_0_72133, HIEFFPLA_NET_0_72134, 
        HIEFFPLA_NET_0_72135, HIEFFPLA_NET_0_72136, 
        HIEFFPLA_NET_0_72137, HIEFFPLA_NET_0_72138, 
        HIEFFPLA_NET_0_72139, HIEFFPLA_NET_0_72140, 
        HIEFFPLA_NET_0_72141, HIEFFPLA_NET_0_72142, 
        HIEFFPLA_NET_0_72143, HIEFFPLA_NET_0_72144, 
        HIEFFPLA_NET_0_72145, HIEFFPLA_NET_0_72146, 
        HIEFFPLA_NET_0_72147, HIEFFPLA_NET_0_72148, 
        HIEFFPLA_NET_0_72149, HIEFFPLA_NET_0_72150, 
        HIEFFPLA_NET_0_72151, HIEFFPLA_NET_0_72152, 
        HIEFFPLA_NET_0_72153, HIEFFPLA_NET_0_72154, 
        HIEFFPLA_NET_0_72155, HIEFFPLA_NET_0_72156, 
        HIEFFPLA_NET_0_72157, HIEFFPLA_NET_0_72158, 
        HIEFFPLA_NET_0_72159, HIEFFPLA_NET_0_72160, 
        HIEFFPLA_NET_0_72161, HIEFFPLA_NET_0_72162, 
        HIEFFPLA_NET_0_72172, HIEFFPLA_NET_0_72173, 
        HIEFFPLA_NET_0_72174, HIEFFPLA_NET_0_72175, 
        HIEFFPLA_NET_0_72176, HIEFFPLA_NET_0_72177, 
        HIEFFPLA_NET_0_72178, HIEFFPLA_NET_0_72179, 
        HIEFFPLA_NET_0_72180, HIEFFPLA_NET_0_72181, 
        HIEFFPLA_NET_0_72182, HIEFFPLA_NET_0_72183, 
        HIEFFPLA_NET_0_72184, HIEFFPLA_NET_0_72185, 
        HIEFFPLA_NET_0_72186, HIEFFPLA_NET_0_72187, 
        HIEFFPLA_NET_0_72188, HIEFFPLA_NET_0_72189, 
        HIEFFPLA_NET_0_72190, HIEFFPLA_NET_0_72191, 
        HIEFFPLA_NET_0_72192, HIEFFPLA_NET_0_72193, 
        HIEFFPLA_NET_0_72194, HIEFFPLA_NET_0_72195, 
        HIEFFPLA_NET_0_72196, HIEFFPLA_NET_0_72197, 
        HIEFFPLA_NET_0_72198, HIEFFPLA_NET_0_72199, 
        HIEFFPLA_NET_0_72200, HIEFFPLA_NET_0_72201, 
        HIEFFPLA_NET_0_72202, HIEFFPLA_NET_0_72203, 
        HIEFFPLA_NET_0_72204, HIEFFPLA_NET_0_72205, 
        HIEFFPLA_NET_0_72206, HIEFFPLA_NET_0_72207, 
        HIEFFPLA_NET_0_72208, HIEFFPLA_NET_0_72209, 
        HIEFFPLA_NET_0_72210, HIEFFPLA_NET_0_72211, 
        HIEFFPLA_NET_0_72212, HIEFFPLA_NET_0_72213, 
        HIEFFPLA_NET_0_72214, HIEFFPLA_NET_0_72215, 
        HIEFFPLA_NET_0_72216, HIEFFPLA_NET_0_72217, 
        HIEFFPLA_NET_0_72218, HIEFFPLA_NET_0_72219, 
        HIEFFPLA_NET_0_72220, HIEFFPLA_NET_0_72221, 
        HIEFFPLA_NET_0_72222, HIEFFPLA_NET_0_72223, 
        HIEFFPLA_NET_0_72224, HIEFFPLA_NET_0_72225, 
        HIEFFPLA_NET_0_72226, HIEFFPLA_NET_0_72227, 
        HIEFFPLA_NET_0_72228, HIEFFPLA_NET_0_72229, 
        HIEFFPLA_NET_0_72230, HIEFFPLA_NET_0_72231, 
        HIEFFPLA_NET_0_72232, HIEFFPLA_NET_0_72233, 
        HIEFFPLA_NET_0_72234, HIEFFPLA_NET_0_72235, 
        HIEFFPLA_NET_0_72236, HIEFFPLA_NET_0_72237, 
        HIEFFPLA_NET_0_72238, HIEFFPLA_NET_0_72239, 
        HIEFFPLA_NET_0_72240, HIEFFPLA_NET_0_72241, 
        HIEFFPLA_NET_0_72242, HIEFFPLA_NET_0_72243, 
        HIEFFPLA_NET_0_72244, HIEFFPLA_NET_0_72245, 
        HIEFFPLA_NET_0_72246, HIEFFPLA_NET_0_72247, 
        HIEFFPLA_NET_0_72248, HIEFFPLA_NET_0_72249, 
        HIEFFPLA_NET_0_72250, HIEFFPLA_NET_0_72251, 
        HIEFFPLA_NET_0_72252, HIEFFPLA_NET_0_72253, 
        HIEFFPLA_NET_0_72254, HIEFFPLA_NET_0_72255, 
        HIEFFPLA_NET_0_72256, HIEFFPLA_NET_0_72257, 
        HIEFFPLA_NET_0_72258, HIEFFPLA_NET_0_72259, 
        HIEFFPLA_NET_0_72260, HIEFFPLA_NET_0_72261, 
        HIEFFPLA_NET_0_72262, HIEFFPLA_NET_0_72263, 
        HIEFFPLA_NET_0_72264, HIEFFPLA_NET_0_72265, 
        HIEFFPLA_NET_0_72266, HIEFFPLA_NET_0_72267, 
        HIEFFPLA_NET_0_72268, HIEFFPLA_NET_0_72269, 
        HIEFFPLA_NET_0_72270, HIEFFPLA_NET_0_72271, 
        HIEFFPLA_NET_0_72272, HIEFFPLA_NET_0_72273, 
        HIEFFPLA_NET_0_72274, HIEFFPLA_NET_0_72275, 
        HIEFFPLA_NET_0_72276, HIEFFPLA_NET_0_72277, 
        HIEFFPLA_NET_0_72278, HIEFFPLA_NET_0_72279, 
        HIEFFPLA_NET_0_72280, HIEFFPLA_NET_0_72281, 
        HIEFFPLA_NET_0_72282, HIEFFPLA_NET_0_72283, 
        HIEFFPLA_NET_0_72284, HIEFFPLA_NET_0_72285, 
        HIEFFPLA_NET_0_72286, HIEFFPLA_NET_0_72287, 
        HIEFFPLA_NET_0_72288, HIEFFPLA_NET_0_72289, 
        HIEFFPLA_NET_0_72290, HIEFFPLA_NET_0_72291, 
        HIEFFPLA_NET_0_72292, HIEFFPLA_NET_0_72293, 
        HIEFFPLA_NET_0_72294, HIEFFPLA_NET_0_72295, 
        HIEFFPLA_NET_0_72296, HIEFFPLA_NET_0_72297, 
        HIEFFPLA_NET_0_72298, HIEFFPLA_NET_0_72299, 
        HIEFFPLA_NET_0_72300, HIEFFPLA_NET_0_72301, 
        HIEFFPLA_NET_0_72302, HIEFFPLA_NET_0_72303, 
        HIEFFPLA_NET_0_72304, HIEFFPLA_NET_0_72305, 
        HIEFFPLA_NET_0_72306, HIEFFPLA_NET_0_72307, 
        HIEFFPLA_NET_0_72308, HIEFFPLA_NET_0_72309, 
        HIEFFPLA_NET_0_72310, HIEFFPLA_NET_0_72311, 
        HIEFFPLA_NET_0_72312, HIEFFPLA_NET_0_72313, 
        HIEFFPLA_NET_0_72314, HIEFFPLA_NET_0_72315, 
        HIEFFPLA_NET_0_72316, HIEFFPLA_NET_0_72317, 
        HIEFFPLA_NET_0_72318, HIEFFPLA_NET_0_72319, 
        HIEFFPLA_NET_0_72320, HIEFFPLA_NET_0_72321, 
        HIEFFPLA_NET_0_72322, HIEFFPLA_NET_0_72323, 
        HIEFFPLA_NET_0_72324, HIEFFPLA_NET_0_72325, 
        HIEFFPLA_NET_0_72326, HIEFFPLA_NET_0_72327, 
        HIEFFPLA_NET_0_72328, HIEFFPLA_NET_0_72329, 
        HIEFFPLA_NET_0_72330, HIEFFPLA_NET_0_72331, 
        HIEFFPLA_NET_0_72332, HIEFFPLA_NET_0_72333, 
        HIEFFPLA_NET_0_72334, HIEFFPLA_NET_0_72335, 
        HIEFFPLA_NET_0_72336, HIEFFPLA_NET_0_72337, 
        HIEFFPLA_NET_0_72338, HIEFFPLA_NET_0_72339, 
        HIEFFPLA_NET_0_72340, HIEFFPLA_NET_0_72341, 
        HIEFFPLA_NET_0_72342, HIEFFPLA_NET_0_72343, 
        HIEFFPLA_NET_0_72344, HIEFFPLA_NET_0_72345, 
        HIEFFPLA_NET_0_72346, HIEFFPLA_NET_0_72347, 
        HIEFFPLA_NET_0_72348, HIEFFPLA_NET_0_72349, 
        HIEFFPLA_NET_0_72350, HIEFFPLA_NET_0_72351, 
        HIEFFPLA_NET_0_72352, HIEFFPLA_NET_0_72353, 
        HIEFFPLA_NET_0_72354, HIEFFPLA_NET_0_72355, 
        HIEFFPLA_NET_0_72356, HIEFFPLA_NET_0_72357, 
        HIEFFPLA_NET_0_72358, HIEFFPLA_NET_0_72359, 
        HIEFFPLA_NET_0_72360, HIEFFPLA_NET_0_72361, 
        HIEFFPLA_NET_0_72362, HIEFFPLA_NET_0_72364, 
        HIEFFPLA_NET_0_72365, HIEFFPLA_NET_0_72366, 
        HIEFFPLA_NET_0_72367, HIEFFPLA_NET_0_72368, 
        HIEFFPLA_NET_0_72369, HIEFFPLA_NET_0_72370, 
        HIEFFPLA_NET_0_72371, HIEFFPLA_NET_0_72372, 
        HIEFFPLA_NET_0_72373, HIEFFPLA_NET_0_72374, 
        HIEFFPLA_NET_0_72375, HIEFFPLA_NET_0_72376, 
        HIEFFPLA_NET_0_72377, HIEFFPLA_NET_0_72378, 
        HIEFFPLA_NET_0_72379, HIEFFPLA_NET_0_72380, 
        HIEFFPLA_NET_0_72381, HIEFFPLA_NET_0_72382, 
        HIEFFPLA_NET_0_72383, HIEFFPLA_NET_0_72384, 
        HIEFFPLA_NET_0_72385, HIEFFPLA_NET_0_72386, 
        HIEFFPLA_NET_0_72387, HIEFFPLA_NET_0_72388, 
        HIEFFPLA_NET_0_72389, HIEFFPLA_NET_0_72390, 
        HIEFFPLA_NET_0_72391, HIEFFPLA_NET_0_72392, 
        HIEFFPLA_NET_0_72393, HIEFFPLA_NET_0_72394, 
        HIEFFPLA_NET_0_72395, HIEFFPLA_NET_0_72396, 
        HIEFFPLA_NET_0_72397, HIEFFPLA_NET_0_72398, 
        HIEFFPLA_NET_0_72399, HIEFFPLA_NET_0_72400, 
        HIEFFPLA_NET_0_72401, HIEFFPLA_NET_0_72402, 
        HIEFFPLA_NET_0_72403, HIEFFPLA_NET_0_72404, 
        HIEFFPLA_NET_0_72405, HIEFFPLA_NET_0_72406, 
        HIEFFPLA_NET_0_72407, HIEFFPLA_NET_0_72408, 
        HIEFFPLA_NET_0_72409, HIEFFPLA_NET_0_72410, 
        HIEFFPLA_NET_0_72411, HIEFFPLA_NET_0_72412, 
        HIEFFPLA_NET_0_72413, HIEFFPLA_NET_0_72414, 
        HIEFFPLA_NET_0_72415, HIEFFPLA_NET_0_72416, 
        HIEFFPLA_NET_0_72417, HIEFFPLA_NET_0_72418, 
        HIEFFPLA_NET_0_72419, HIEFFPLA_NET_0_72420, 
        HIEFFPLA_NET_0_72421, HIEFFPLA_NET_0_72422, 
        HIEFFPLA_NET_0_72423, HIEFFPLA_NET_0_72424, 
        HIEFFPLA_NET_0_72425, HIEFFPLA_NET_0_72426, 
        HIEFFPLA_NET_0_72427, HIEFFPLA_NET_0_72428, 
        HIEFFPLA_NET_0_72429, HIEFFPLA_NET_0_72430, 
        HIEFFPLA_NET_0_72431, HIEFFPLA_NET_0_72432, 
        HIEFFPLA_NET_0_72433, HIEFFPLA_NET_0_72434, 
        HIEFFPLA_NET_0_72435, HIEFFPLA_NET_0_72436, 
        HIEFFPLA_NET_0_72437, HIEFFPLA_NET_0_72438, 
        HIEFFPLA_NET_0_72439, HIEFFPLA_NET_0_72440, 
        HIEFFPLA_NET_0_72441, HIEFFPLA_NET_0_72442, 
        HIEFFPLA_NET_0_72443, HIEFFPLA_NET_0_72444, 
        HIEFFPLA_NET_0_72445, HIEFFPLA_NET_0_72446, 
        HIEFFPLA_NET_0_72447, HIEFFPLA_NET_0_72448, 
        HIEFFPLA_NET_0_72449, HIEFFPLA_NET_0_72450, 
        HIEFFPLA_NET_0_72451, HIEFFPLA_NET_0_72452, 
        HIEFFPLA_NET_0_72453, HIEFFPLA_NET_0_72454, 
        HIEFFPLA_NET_0_72455, HIEFFPLA_NET_0_72456, 
        HIEFFPLA_NET_0_72457, HIEFFPLA_NET_0_72458, 
        HIEFFPLA_NET_0_72459, HIEFFPLA_NET_0_72460, 
        HIEFFPLA_NET_0_72461, HIEFFPLA_NET_0_72462, 
        HIEFFPLA_NET_0_72463, HIEFFPLA_NET_0_72464, 
        HIEFFPLA_NET_0_72465, HIEFFPLA_NET_0_72466, 
        HIEFFPLA_NET_0_72467, HIEFFPLA_NET_0_72468, 
        HIEFFPLA_NET_0_72469, HIEFFPLA_NET_0_72470, 
        HIEFFPLA_NET_0_72471, HIEFFPLA_NET_0_72472, 
        HIEFFPLA_NET_0_72473, HIEFFPLA_NET_0_72474, 
        HIEFFPLA_NET_0_72475, HIEFFPLA_NET_0_72476, 
        HIEFFPLA_NET_0_72477, HIEFFPLA_NET_0_72478, 
        HIEFFPLA_NET_0_72479, HIEFFPLA_NET_0_72480, 
        HIEFFPLA_NET_0_72481, HIEFFPLA_NET_0_72482, 
        HIEFFPLA_NET_0_72483, HIEFFPLA_NET_0_72484, 
        HIEFFPLA_NET_0_72485, HIEFFPLA_NET_0_72486, 
        HIEFFPLA_NET_0_72487, HIEFFPLA_NET_0_72488, 
        HIEFFPLA_NET_0_72489, HIEFFPLA_NET_0_72490, 
        HIEFFPLA_NET_0_72491, HIEFFPLA_NET_0_72492, 
        HIEFFPLA_NET_0_72493, HIEFFPLA_NET_0_72494, 
        HIEFFPLA_NET_0_72495, HIEFFPLA_NET_0_72496, 
        HIEFFPLA_NET_0_72497, HIEFFPLA_NET_0_72498, 
        HIEFFPLA_NET_0_72499, HIEFFPLA_NET_0_72500, 
        HIEFFPLA_NET_0_72501, HIEFFPLA_NET_0_72502, 
        HIEFFPLA_NET_0_72503, HIEFFPLA_NET_0_72504, 
        HIEFFPLA_NET_0_72505, HIEFFPLA_NET_0_72506, 
        HIEFFPLA_NET_0_72507, HIEFFPLA_NET_0_72508, 
        HIEFFPLA_NET_0_72509, HIEFFPLA_NET_0_72510, 
        HIEFFPLA_NET_0_72511, HIEFFPLA_NET_0_72512, 
        HIEFFPLA_NET_0_72513, HIEFFPLA_NET_0_72514, 
        HIEFFPLA_NET_0_72515, HIEFFPLA_NET_0_72516, 
        HIEFFPLA_NET_0_72517, HIEFFPLA_NET_0_72518, 
        HIEFFPLA_NET_0_72519, HIEFFPLA_NET_0_72520, 
        HIEFFPLA_NET_0_72521, HIEFFPLA_NET_0_72522, 
        HIEFFPLA_NET_0_72523, HIEFFPLA_NET_0_72524, 
        HIEFFPLA_NET_0_72525, HIEFFPLA_NET_0_72526, 
        HIEFFPLA_NET_0_72527, HIEFFPLA_NET_0_72528, 
        HIEFFPLA_NET_0_72529, HIEFFPLA_NET_0_72530, 
        HIEFFPLA_NET_0_72531, HIEFFPLA_NET_0_72532, 
        HIEFFPLA_NET_0_72533, HIEFFPLA_NET_0_72534, 
        HIEFFPLA_NET_0_72535, HIEFFPLA_NET_0_72536, 
        HIEFFPLA_NET_0_72537, HIEFFPLA_NET_0_72538, 
        HIEFFPLA_NET_0_72539, HIEFFPLA_NET_0_72540, 
        HIEFFPLA_NET_0_72541, HIEFFPLA_NET_0_72542, 
        HIEFFPLA_NET_0_72543, HIEFFPLA_NET_0_72544, 
        HIEFFPLA_NET_0_72545, HIEFFPLA_NET_0_72546, 
        HIEFFPLA_NET_0_72547, HIEFFPLA_NET_0_72548, 
        HIEFFPLA_NET_0_72549, HIEFFPLA_NET_0_72550, 
        HIEFFPLA_NET_0_72551, HIEFFPLA_NET_0_72552, 
        HIEFFPLA_NET_0_72553, HIEFFPLA_NET_0_72554, 
        HIEFFPLA_NET_0_72555, HIEFFPLA_NET_0_72556, 
        HIEFFPLA_NET_0_72557, HIEFFPLA_NET_0_72558, 
        HIEFFPLA_NET_0_72559, HIEFFPLA_NET_0_72560, 
        HIEFFPLA_NET_0_72561, HIEFFPLA_NET_0_72562, 
        HIEFFPLA_NET_0_72563, HIEFFPLA_NET_0_72564, 
        HIEFFPLA_NET_0_72565, HIEFFPLA_NET_0_72566, 
        HIEFFPLA_NET_0_72567, HIEFFPLA_NET_0_72568, 
        HIEFFPLA_NET_0_72569, HIEFFPLA_NET_0_72570, 
        HIEFFPLA_NET_0_72571, HIEFFPLA_NET_0_72572, 
        HIEFFPLA_NET_0_72573, HIEFFPLA_NET_0_72574, 
        HIEFFPLA_NET_0_72575, HIEFFPLA_NET_0_72576, 
        HIEFFPLA_NET_0_72577, HIEFFPLA_NET_0_72578, 
        HIEFFPLA_NET_0_72579, HIEFFPLA_NET_0_72580, 
        HIEFFPLA_NET_0_72581, HIEFFPLA_NET_0_72582, 
        HIEFFPLA_NET_0_72583, HIEFFPLA_NET_0_72584, 
        HIEFFPLA_NET_0_72585, HIEFFPLA_NET_0_72586, 
        HIEFFPLA_NET_0_72587, HIEFFPLA_NET_0_72588, 
        HIEFFPLA_NET_0_72589, HIEFFPLA_NET_0_72590, 
        HIEFFPLA_NET_0_72591, HIEFFPLA_NET_0_72592, 
        HIEFFPLA_NET_0_72593, HIEFFPLA_NET_0_72594, 
        HIEFFPLA_NET_0_72595, HIEFFPLA_NET_0_72596, 
        HIEFFPLA_NET_0_72597, HIEFFPLA_NET_0_72598, 
        HIEFFPLA_NET_0_72599, HIEFFPLA_NET_0_72600, 
        HIEFFPLA_NET_0_72601, HIEFFPLA_NET_0_72602, 
        HIEFFPLA_NET_0_72603, HIEFFPLA_NET_0_72604, 
        HIEFFPLA_NET_0_72605, HIEFFPLA_NET_0_72606, 
        HIEFFPLA_NET_0_72607, HIEFFPLA_NET_0_72608, 
        HIEFFPLA_NET_0_72609, HIEFFPLA_NET_0_72610, 
        HIEFFPLA_NET_0_72611, HIEFFPLA_NET_0_72612, 
        HIEFFPLA_NET_0_72613, HIEFFPLA_NET_0_72614, 
        HIEFFPLA_NET_0_72615, HIEFFPLA_NET_0_72616, 
        HIEFFPLA_NET_0_72617, HIEFFPLA_NET_0_72618, 
        HIEFFPLA_NET_0_72619, HIEFFPLA_NET_0_72620, 
        HIEFFPLA_NET_0_72621, HIEFFPLA_NET_0_72622, 
        HIEFFPLA_NET_0_72623, HIEFFPLA_NET_0_72624, 
        HIEFFPLA_NET_0_72625, HIEFFPLA_NET_0_72626, 
        HIEFFPLA_NET_0_72627, HIEFFPLA_NET_0_72628, 
        HIEFFPLA_NET_0_72629, HIEFFPLA_NET_0_72630, 
        HIEFFPLA_NET_0_72631, HIEFFPLA_NET_0_72632, 
        HIEFFPLA_NET_0_72633, HIEFFPLA_NET_0_72634, 
        HIEFFPLA_NET_0_72635, HIEFFPLA_NET_0_72636, 
        HIEFFPLA_NET_0_72637, HIEFFPLA_NET_0_72638, 
        HIEFFPLA_NET_0_72639, HIEFFPLA_NET_0_72640, 
        HIEFFPLA_NET_0_72641, HIEFFPLA_NET_0_72642, 
        HIEFFPLA_NET_0_72643, HIEFFPLA_NET_0_72645, 
        HIEFFPLA_NET_0_72646, HIEFFPLA_NET_0_72647, 
        HIEFFPLA_NET_0_72648, HIEFFPLA_NET_0_72649, 
        HIEFFPLA_NET_0_72650, HIEFFPLA_NET_0_72651, 
        HIEFFPLA_NET_0_72652, HIEFFPLA_NET_0_72653, 
        HIEFFPLA_NET_0_72654, HIEFFPLA_NET_0_72655, 
        HIEFFPLA_NET_0_72656, HIEFFPLA_NET_0_72657, 
        HIEFFPLA_NET_0_72658, HIEFFPLA_NET_0_72659, 
        HIEFFPLA_NET_0_72660, HIEFFPLA_NET_0_72661, 
        HIEFFPLA_NET_0_72662, HIEFFPLA_NET_0_72663, 
        HIEFFPLA_NET_0_72664, HIEFFPLA_NET_0_72665, 
        HIEFFPLA_NET_0_72666, HIEFFPLA_NET_0_72667, 
        HIEFFPLA_NET_0_72668, HIEFFPLA_NET_0_72669, 
        HIEFFPLA_NET_0_72670, HIEFFPLA_NET_0_72671, 
        HIEFFPLA_NET_0_72672, HIEFFPLA_NET_0_72673, 
        HIEFFPLA_NET_0_72674, HIEFFPLA_NET_0_72675, 
        HIEFFPLA_NET_0_72676, HIEFFPLA_NET_0_72677, 
        HIEFFPLA_NET_0_72678, HIEFFPLA_NET_0_72679, 
        HIEFFPLA_NET_0_72680, HIEFFPLA_NET_0_72681, 
        HIEFFPLA_NET_0_72682, HIEFFPLA_NET_0_72683, 
        HIEFFPLA_NET_0_72684, HIEFFPLA_NET_0_72685, 
        HIEFFPLA_NET_0_72686, HIEFFPLA_NET_0_72687, 
        HIEFFPLA_NET_0_72688, HIEFFPLA_NET_0_72689, 
        HIEFFPLA_NET_0_72690, HIEFFPLA_NET_0_72691, 
        HIEFFPLA_NET_0_72692, HIEFFPLA_NET_0_72693, 
        HIEFFPLA_NET_0_72694, HIEFFPLA_NET_0_72695, 
        HIEFFPLA_NET_0_72696, HIEFFPLA_NET_0_72697, 
        HIEFFPLA_NET_0_72698, HIEFFPLA_NET_0_72699, 
        HIEFFPLA_NET_0_72700, HIEFFPLA_NET_0_72701, 
        HIEFFPLA_NET_0_72702, HIEFFPLA_NET_0_72703, 
        HIEFFPLA_NET_0_72704, HIEFFPLA_NET_0_72705, 
        HIEFFPLA_NET_0_72706, HIEFFPLA_NET_0_72707, 
        HIEFFPLA_NET_0_72708, HIEFFPLA_NET_0_72709, 
        HIEFFPLA_NET_0_72710, HIEFFPLA_NET_0_72711, 
        HIEFFPLA_NET_0_72712, HIEFFPLA_NET_0_72713, 
        HIEFFPLA_NET_0_72714, HIEFFPLA_NET_0_72715, 
        HIEFFPLA_NET_0_72716, HIEFFPLA_NET_0_72717, 
        HIEFFPLA_NET_0_72718, HIEFFPLA_NET_0_72719, 
        HIEFFPLA_NET_0_72720, HIEFFPLA_NET_0_72721, 
        HIEFFPLA_NET_0_72722, HIEFFPLA_NET_0_72723, 
        HIEFFPLA_NET_0_72724, HIEFFPLA_NET_0_72725, 
        HIEFFPLA_NET_0_72726, HIEFFPLA_NET_0_72727, 
        HIEFFPLA_NET_0_72728, HIEFFPLA_NET_0_72729, 
        HIEFFPLA_NET_0_72730, HIEFFPLA_NET_0_72731, 
        HIEFFPLA_NET_0_72732, HIEFFPLA_NET_0_72733, 
        HIEFFPLA_NET_0_72734, HIEFFPLA_NET_0_72735, 
        HIEFFPLA_NET_0_72736, HIEFFPLA_NET_0_72737, 
        HIEFFPLA_NET_0_72738, HIEFFPLA_NET_0_72739, 
        HIEFFPLA_NET_0_72740, HIEFFPLA_NET_0_72741, 
        HIEFFPLA_NET_0_72742, HIEFFPLA_NET_0_72743, 
        HIEFFPLA_NET_0_72744, HIEFFPLA_NET_0_72745, 
        HIEFFPLA_NET_0_72746, HIEFFPLA_NET_0_72747, 
        HIEFFPLA_NET_0_72748, HIEFFPLA_NET_0_72749, 
        HIEFFPLA_NET_0_72750, HIEFFPLA_NET_0_72751, 
        HIEFFPLA_NET_0_72752, HIEFFPLA_NET_0_72753, 
        HIEFFPLA_NET_0_72754, HIEFFPLA_NET_0_72755, 
        HIEFFPLA_NET_0_72756, HIEFFPLA_NET_0_72757, 
        HIEFFPLA_NET_0_72758, HIEFFPLA_NET_0_72759, 
        HIEFFPLA_NET_0_72760, HIEFFPLA_NET_0_72761, 
        HIEFFPLA_NET_0_72762, HIEFFPLA_NET_0_72763, 
        HIEFFPLA_NET_0_72764, HIEFFPLA_NET_0_72765, 
        HIEFFPLA_NET_0_72766, HIEFFPLA_NET_0_72767, 
        HIEFFPLA_NET_0_72768, HIEFFPLA_NET_0_72769, 
        HIEFFPLA_NET_0_72770, HIEFFPLA_NET_0_72771, 
        HIEFFPLA_NET_0_72772, HIEFFPLA_NET_0_72773, 
        HIEFFPLA_NET_0_72774, HIEFFPLA_NET_0_72775, 
        HIEFFPLA_NET_0_72776, HIEFFPLA_NET_0_72777, 
        HIEFFPLA_NET_0_72778, HIEFFPLA_NET_0_72779, 
        HIEFFPLA_NET_0_72780, HIEFFPLA_NET_0_72781, 
        HIEFFPLA_NET_0_72782, HIEFFPLA_NET_0_72783, 
        HIEFFPLA_NET_0_72784, HIEFFPLA_NET_0_72785, 
        HIEFFPLA_NET_0_72786, HIEFFPLA_NET_0_72787, 
        HIEFFPLA_NET_0_72788, HIEFFPLA_NET_0_72789, 
        HIEFFPLA_NET_0_72790, HIEFFPLA_NET_0_72791, 
        HIEFFPLA_NET_0_72792, HIEFFPLA_NET_0_72793, 
        HIEFFPLA_NET_0_72794, HIEFFPLA_NET_0_72795, 
        HIEFFPLA_NET_0_72796, HIEFFPLA_NET_0_72797, 
        HIEFFPLA_NET_0_72798, HIEFFPLA_NET_0_72799, 
        HIEFFPLA_NET_0_72800, HIEFFPLA_NET_0_72801, 
        HIEFFPLA_NET_0_72802, HIEFFPLA_NET_0_72803, 
        HIEFFPLA_NET_0_72804, HIEFFPLA_NET_0_72805, 
        HIEFFPLA_NET_0_72806, HIEFFPLA_NET_0_72807, 
        HIEFFPLA_NET_0_72808, HIEFFPLA_NET_0_72809, 
        HIEFFPLA_NET_0_72810, HIEFFPLA_NET_0_72811, 
        HIEFFPLA_NET_0_72812, HIEFFPLA_NET_0_72813, 
        HIEFFPLA_NET_0_72814, HIEFFPLA_NET_0_72815, 
        HIEFFPLA_NET_0_72816, HIEFFPLA_NET_0_72817, 
        HIEFFPLA_NET_0_72818, HIEFFPLA_NET_0_72819, 
        HIEFFPLA_NET_0_72820, HIEFFPLA_NET_0_72821, 
        HIEFFPLA_NET_0_72822, HIEFFPLA_NET_0_72823, 
        HIEFFPLA_NET_0_72824, HIEFFPLA_NET_0_72825, 
        HIEFFPLA_NET_0_72826, HIEFFPLA_NET_0_72827, 
        HIEFFPLA_NET_0_72828, HIEFFPLA_NET_0_72829, 
        HIEFFPLA_NET_0_72830, HIEFFPLA_NET_0_72831, 
        HIEFFPLA_NET_0_72832, HIEFFPLA_NET_0_72833, 
        HIEFFPLA_NET_0_72834, HIEFFPLA_NET_0_72835, 
        HIEFFPLA_NET_0_72836, HIEFFPLA_NET_0_72837, 
        HIEFFPLA_NET_0_72838, HIEFFPLA_NET_0_72839, 
        HIEFFPLA_NET_0_72840, HIEFFPLA_NET_0_72841, 
        HIEFFPLA_NET_0_72842, HIEFFPLA_NET_0_72843, 
        HIEFFPLA_NET_0_72844, HIEFFPLA_NET_0_72845, 
        HIEFFPLA_NET_0_72846, HIEFFPLA_NET_0_72847, 
        HIEFFPLA_NET_0_72848, HIEFFPLA_NET_0_72849, 
        HIEFFPLA_NET_0_72850, HIEFFPLA_NET_0_72851, 
        HIEFFPLA_NET_0_72852, HIEFFPLA_NET_0_72853, 
        HIEFFPLA_NET_0_72854, HIEFFPLA_NET_0_72855, 
        HIEFFPLA_NET_0_72856, HIEFFPLA_NET_0_72857, 
        HIEFFPLA_NET_0_72858, HIEFFPLA_NET_0_72859, 
        HIEFFPLA_NET_0_72860, HIEFFPLA_NET_0_72861, 
        HIEFFPLA_NET_0_72862, HIEFFPLA_NET_0_72863, 
        HIEFFPLA_NET_0_72864, HIEFFPLA_NET_0_72865, 
        HIEFFPLA_NET_0_72866, HIEFFPLA_NET_0_72867, 
        HIEFFPLA_NET_0_72868, HIEFFPLA_NET_0_72869, 
        HIEFFPLA_NET_0_72870, HIEFFPLA_NET_0_72871, 
        HIEFFPLA_NET_0_72872, HIEFFPLA_NET_0_72873, 
        HIEFFPLA_NET_0_72874, HIEFFPLA_NET_0_72875, 
        HIEFFPLA_NET_0_72876, HIEFFPLA_NET_0_72877, 
        HIEFFPLA_NET_0_72878, HIEFFPLA_NET_0_72879, 
        HIEFFPLA_NET_0_72880, HIEFFPLA_NET_0_72881, 
        HIEFFPLA_NET_0_72882, HIEFFPLA_NET_0_72883, 
        HIEFFPLA_NET_0_72884, HIEFFPLA_NET_0_72885, 
        HIEFFPLA_NET_0_72886, HIEFFPLA_NET_0_72887, 
        HIEFFPLA_NET_0_72888, HIEFFPLA_NET_0_72889, 
        HIEFFPLA_NET_0_72890, HIEFFPLA_NET_0_72891, 
        HIEFFPLA_NET_0_72892, HIEFFPLA_NET_0_72893, 
        HIEFFPLA_NET_0_72894, HIEFFPLA_NET_0_72895, 
        HIEFFPLA_NET_0_72896, HIEFFPLA_NET_0_72897, 
        HIEFFPLA_NET_0_72898, HIEFFPLA_NET_0_72899, 
        HIEFFPLA_NET_0_72900, HIEFFPLA_NET_0_72901, 
        HIEFFPLA_NET_0_72902, HIEFFPLA_NET_0_72903, 
        HIEFFPLA_NET_0_72904, HIEFFPLA_NET_0_72905, 
        HIEFFPLA_NET_0_72906, HIEFFPLA_NET_0_72907, 
        HIEFFPLA_NET_0_72908, HIEFFPLA_NET_0_72909, 
        HIEFFPLA_NET_0_72910, HIEFFPLA_NET_0_72911, 
        HIEFFPLA_NET_0_72912, HIEFFPLA_NET_0_72913, 
        HIEFFPLA_NET_0_72914, HIEFFPLA_NET_0_72915, 
        HIEFFPLA_NET_0_72916, HIEFFPLA_NET_0_72917, 
        HIEFFPLA_NET_0_72918, HIEFFPLA_NET_0_72919, 
        HIEFFPLA_NET_0_72920, HIEFFPLA_NET_0_72921, 
        HIEFFPLA_NET_0_72922, HIEFFPLA_NET_0_72923, 
        HIEFFPLA_NET_0_72924, HIEFFPLA_NET_0_72925, 
        HIEFFPLA_NET_0_72926, HIEFFPLA_NET_0_72927, 
        HIEFFPLA_NET_0_72928, HIEFFPLA_NET_0_72929, 
        HIEFFPLA_NET_0_72930, HIEFFPLA_NET_0_72931, 
        HIEFFPLA_NET_0_72932, HIEFFPLA_NET_0_72933, 
        HIEFFPLA_NET_0_72934, HIEFFPLA_NET_0_72935, 
        HIEFFPLA_NET_0_72936, HIEFFPLA_NET_0_72937, 
        HIEFFPLA_NET_0_72938, HIEFFPLA_NET_0_72939, 
        HIEFFPLA_NET_0_72940, HIEFFPLA_NET_0_72941, 
        HIEFFPLA_NET_0_72942, HIEFFPLA_NET_0_72943, 
        HIEFFPLA_NET_0_72944, HIEFFPLA_NET_0_72945, 
        HIEFFPLA_NET_0_72946, HIEFFPLA_NET_0_72947, 
        HIEFFPLA_NET_0_72948, HIEFFPLA_NET_0_72949, 
        HIEFFPLA_NET_0_72950, HIEFFPLA_NET_0_72951, 
        HIEFFPLA_NET_0_72952, HIEFFPLA_NET_0_72953, 
        HIEFFPLA_NET_0_72954, HIEFFPLA_NET_0_72955, 
        HIEFFPLA_NET_0_72956, HIEFFPLA_NET_0_72957, 
        HIEFFPLA_NET_0_72958, HIEFFPLA_NET_0_72959, 
        HIEFFPLA_NET_0_72960, HIEFFPLA_NET_0_72961, 
        HIEFFPLA_NET_0_72962, HIEFFPLA_NET_0_72963, 
        HIEFFPLA_NET_0_72964, HIEFFPLA_NET_0_72965, 
        HIEFFPLA_NET_0_72966, HIEFFPLA_NET_0_72967, 
        HIEFFPLA_NET_0_72968, HIEFFPLA_NET_0_72969, 
        HIEFFPLA_NET_0_72970, HIEFFPLA_NET_0_72971, 
        HIEFFPLA_NET_0_72972, HIEFFPLA_NET_0_72973, 
        HIEFFPLA_NET_0_72974, HIEFFPLA_NET_0_72975, 
        HIEFFPLA_NET_0_72976, HIEFFPLA_NET_0_72977, 
        HIEFFPLA_NET_0_72978, HIEFFPLA_NET_0_72979, 
        HIEFFPLA_NET_0_72980, HIEFFPLA_NET_0_72981, 
        HIEFFPLA_NET_0_72982, HIEFFPLA_NET_0_72983, 
        HIEFFPLA_NET_0_72984, HIEFFPLA_NET_0_72985, 
        HIEFFPLA_NET_0_72986, HIEFFPLA_NET_0_72987, 
        HIEFFPLA_NET_0_72988, HIEFFPLA_NET_0_72989, 
        HIEFFPLA_NET_0_72990, HIEFFPLA_NET_0_72991, 
        HIEFFPLA_NET_0_72992, HIEFFPLA_NET_0_72993, 
        HIEFFPLA_NET_0_72994, HIEFFPLA_NET_0_72995, 
        HIEFFPLA_NET_0_72996, HIEFFPLA_NET_0_72997, 
        HIEFFPLA_NET_0_72998, HIEFFPLA_NET_0_72999, 
        HIEFFPLA_NET_0_73000, HIEFFPLA_NET_0_73001, 
        HIEFFPLA_NET_0_73002, HIEFFPLA_NET_0_73003, 
        HIEFFPLA_NET_0_73004, HIEFFPLA_NET_0_73005, 
        HIEFFPLA_NET_0_73006, HIEFFPLA_NET_0_73007, 
        HIEFFPLA_NET_0_73008, HIEFFPLA_NET_0_73009, 
        HIEFFPLA_NET_0_73010, HIEFFPLA_NET_0_73011, 
        HIEFFPLA_NET_0_73012, HIEFFPLA_NET_0_73013, 
        HIEFFPLA_NET_0_73014, HIEFFPLA_NET_0_73015, 
        HIEFFPLA_NET_0_73016, HIEFFPLA_NET_0_73017, 
        HIEFFPLA_NET_0_73018, HIEFFPLA_NET_0_73019, 
        HIEFFPLA_NET_0_73020, HIEFFPLA_NET_0_73021, 
        HIEFFPLA_NET_0_73022, HIEFFPLA_NET_0_73023, 
        HIEFFPLA_NET_0_73024, HIEFFPLA_NET_0_73025, 
        HIEFFPLA_NET_0_73026, HIEFFPLA_NET_0_73027, 
        HIEFFPLA_NET_0_73028, HIEFFPLA_NET_0_73029, 
        HIEFFPLA_NET_0_73030, HIEFFPLA_NET_0_73031, 
        HIEFFPLA_NET_0_73032, HIEFFPLA_NET_0_73033, 
        HIEFFPLA_NET_0_73034, HIEFFPLA_NET_0_73035, 
        HIEFFPLA_NET_0_73036, HIEFFPLA_NET_0_73037, 
        HIEFFPLA_NET_0_73038, HIEFFPLA_NET_0_73039, 
        HIEFFPLA_NET_0_73040, HIEFFPLA_NET_0_73041, 
        HIEFFPLA_NET_0_73042, HIEFFPLA_NET_0_73043, 
        HIEFFPLA_NET_0_73044, HIEFFPLA_NET_0_73045, 
        HIEFFPLA_NET_0_73046, HIEFFPLA_NET_0_73047, 
        HIEFFPLA_NET_0_73048, HIEFFPLA_NET_0_73049, 
        HIEFFPLA_NET_0_73050, HIEFFPLA_NET_0_73051, 
        HIEFFPLA_NET_0_73052, HIEFFPLA_NET_0_73053, 
        HIEFFPLA_NET_0_73054, HIEFFPLA_NET_0_73055, 
        HIEFFPLA_NET_0_73056, HIEFFPLA_NET_0_73057, 
        HIEFFPLA_NET_0_73058, HIEFFPLA_NET_0_73059, 
        HIEFFPLA_NET_0_73060, HIEFFPLA_NET_0_73061, 
        HIEFFPLA_NET_0_73062, HIEFFPLA_NET_0_73063, 
        HIEFFPLA_NET_0_73064, HIEFFPLA_NET_0_73065, 
        HIEFFPLA_NET_0_73066, HIEFFPLA_NET_0_73067, 
        HIEFFPLA_NET_0_73068, HIEFFPLA_NET_0_73069, 
        HIEFFPLA_NET_0_73070, HIEFFPLA_NET_0_73071, 
        HIEFFPLA_NET_0_73072, HIEFFPLA_NET_0_73073, 
        HIEFFPLA_NET_0_73075, HIEFFPLA_NET_0_73076, 
        HIEFFPLA_NET_0_73077, HIEFFPLA_NET_0_73078, 
        HIEFFPLA_NET_0_73079, HIEFFPLA_NET_0_73080, 
        HIEFFPLA_NET_0_73081, HIEFFPLA_NET_0_73082, 
        HIEFFPLA_NET_0_73083, HIEFFPLA_NET_0_73084, 
        HIEFFPLA_NET_0_73085, HIEFFPLA_NET_0_73086, 
        HIEFFPLA_NET_0_73087, HIEFFPLA_NET_0_73088, 
        HIEFFPLA_NET_0_73089, HIEFFPLA_NET_0_73090, 
        HIEFFPLA_NET_0_73091, HIEFFPLA_NET_0_73092, 
        HIEFFPLA_NET_0_73093, HIEFFPLA_NET_0_73094, 
        HIEFFPLA_NET_0_73095, HIEFFPLA_NET_0_73096, 
        HIEFFPLA_NET_0_73097, HIEFFPLA_NET_0_73098, 
        HIEFFPLA_NET_0_73099, HIEFFPLA_NET_0_73100, 
        HIEFFPLA_NET_0_73101, HIEFFPLA_NET_0_73102, 
        HIEFFPLA_NET_0_73103, HIEFFPLA_NET_0_73104, 
        HIEFFPLA_NET_0_73105, HIEFFPLA_NET_0_73106, 
        HIEFFPLA_NET_0_73107, HIEFFPLA_NET_0_73108, 
        HIEFFPLA_NET_0_73109, HIEFFPLA_NET_0_73110, 
        HIEFFPLA_NET_0_73111, HIEFFPLA_NET_0_73112, 
        HIEFFPLA_NET_0_73113, HIEFFPLA_NET_0_73114, 
        HIEFFPLA_NET_0_73115, HIEFFPLA_NET_0_73116, 
        HIEFFPLA_NET_0_73117, HIEFFPLA_NET_0_73118, 
        HIEFFPLA_NET_0_73119, HIEFFPLA_NET_0_73120, 
        HIEFFPLA_NET_0_73121, HIEFFPLA_NET_0_73122, 
        HIEFFPLA_NET_0_73123, HIEFFPLA_NET_0_73124, 
        HIEFFPLA_NET_0_73125, HIEFFPLA_NET_0_73126, 
        HIEFFPLA_NET_0_73127, HIEFFPLA_NET_0_73128, 
        HIEFFPLA_NET_0_73129, HIEFFPLA_NET_0_73130, 
        HIEFFPLA_NET_0_73131, HIEFFPLA_NET_0_73132, 
        HIEFFPLA_NET_0_73133, HIEFFPLA_NET_0_73134, 
        HIEFFPLA_NET_0_73135, HIEFFPLA_NET_0_73136, 
        HIEFFPLA_NET_0_73137, HIEFFPLA_NET_0_73138, 
        HIEFFPLA_NET_0_73139, HIEFFPLA_NET_0_73140, 
        HIEFFPLA_NET_0_73141, HIEFFPLA_NET_0_73142, 
        HIEFFPLA_NET_0_73143, HIEFFPLA_NET_0_73144, 
        HIEFFPLA_NET_0_73145, HIEFFPLA_NET_0_73146, 
        HIEFFPLA_NET_0_73147, HIEFFPLA_NET_0_73148, 
        HIEFFPLA_NET_0_73149, HIEFFPLA_NET_0_73150, 
        HIEFFPLA_NET_0_73151, HIEFFPLA_NET_0_73152, 
        HIEFFPLA_NET_0_73153, HIEFFPLA_NET_0_73154, 
        HIEFFPLA_NET_0_73155, HIEFFPLA_NET_0_73156, 
        HIEFFPLA_NET_0_73157, HIEFFPLA_NET_0_73158, 
        HIEFFPLA_NET_0_73159, HIEFFPLA_NET_0_73160, 
        HIEFFPLA_NET_0_73161, HIEFFPLA_NET_0_73162, 
        HIEFFPLA_NET_0_73163, HIEFFPLA_NET_0_73164, 
        HIEFFPLA_NET_0_73165, HIEFFPLA_NET_0_73166, 
        HIEFFPLA_NET_0_73167, HIEFFPLA_NET_0_73168, 
        HIEFFPLA_NET_0_73169, HIEFFPLA_NET_0_73170, 
        HIEFFPLA_NET_0_73171, HIEFFPLA_NET_0_73172, 
        HIEFFPLA_NET_0_73173, HIEFFPLA_NET_0_73174, 
        HIEFFPLA_NET_0_73175, HIEFFPLA_NET_0_73176, 
        HIEFFPLA_NET_0_73177, HIEFFPLA_NET_0_73178, 
        HIEFFPLA_NET_0_73179, HIEFFPLA_NET_0_73180, 
        HIEFFPLA_NET_0_73181, HIEFFPLA_NET_0_73182, 
        HIEFFPLA_NET_0_73183, HIEFFPLA_NET_0_73184, 
        HIEFFPLA_NET_0_73185, HIEFFPLA_NET_0_73186, 
        HIEFFPLA_NET_0_73187, HIEFFPLA_NET_0_73188, 
        HIEFFPLA_NET_0_73189, HIEFFPLA_NET_0_73190, 
        HIEFFPLA_NET_0_73191, HIEFFPLA_NET_0_73192, 
        HIEFFPLA_NET_0_73193, HIEFFPLA_NET_0_73194, 
        HIEFFPLA_NET_0_73195, HIEFFPLA_NET_0_73196, 
        HIEFFPLA_NET_0_73197, HIEFFPLA_NET_0_73198, 
        HIEFFPLA_NET_0_73199, HIEFFPLA_NET_0_73200, 
        HIEFFPLA_NET_0_73201, HIEFFPLA_NET_0_73202, 
        HIEFFPLA_NET_0_73203, HIEFFPLA_NET_0_73204, 
        HIEFFPLA_NET_0_73205, HIEFFPLA_NET_0_73206, 
        HIEFFPLA_NET_0_73207, HIEFFPLA_NET_0_73208, 
        HIEFFPLA_NET_0_73209, HIEFFPLA_NET_0_73210, 
        HIEFFPLA_NET_0_73211, HIEFFPLA_NET_0_73212, 
        HIEFFPLA_NET_0_73213, HIEFFPLA_NET_0_73214, 
        HIEFFPLA_NET_0_73215, HIEFFPLA_NET_0_73216, 
        HIEFFPLA_NET_0_73217, HIEFFPLA_NET_0_73218, 
        HIEFFPLA_NET_0_73219, HIEFFPLA_NET_0_73220, 
        HIEFFPLA_NET_0_73221, HIEFFPLA_NET_0_73222, 
        HIEFFPLA_NET_0_73223, HIEFFPLA_NET_0_73224, 
        HIEFFPLA_NET_0_73225, HIEFFPLA_NET_0_73226, 
        HIEFFPLA_NET_0_73227, HIEFFPLA_NET_0_73228, 
        HIEFFPLA_NET_0_73229, HIEFFPLA_NET_0_73230, 
        HIEFFPLA_NET_0_73231, HIEFFPLA_NET_0_73232, 
        HIEFFPLA_NET_0_73233, HIEFFPLA_NET_0_73234, 
        HIEFFPLA_NET_0_73235, HIEFFPLA_NET_0_73236, 
        HIEFFPLA_NET_0_73237, HIEFFPLA_NET_0_73238, 
        HIEFFPLA_NET_0_73239, HIEFFPLA_NET_0_73240, 
        HIEFFPLA_NET_0_73241, HIEFFPLA_NET_0_73242, 
        HIEFFPLA_NET_0_73243, HIEFFPLA_NET_0_73244, 
        HIEFFPLA_NET_0_73245, HIEFFPLA_NET_0_73246, 
        HIEFFPLA_NET_0_73247, HIEFFPLA_NET_0_73248, 
        HIEFFPLA_NET_0_73249, HIEFFPLA_NET_0_73250, 
        HIEFFPLA_NET_0_73251, HIEFFPLA_NET_0_73252, 
        HIEFFPLA_NET_0_73253, HIEFFPLA_NET_0_73254, 
        HIEFFPLA_NET_0_73255, HIEFFPLA_NET_0_73256, 
        HIEFFPLA_NET_0_73257, HIEFFPLA_NET_0_73258, 
        HIEFFPLA_NET_0_73259, HIEFFPLA_NET_0_73260, 
        HIEFFPLA_NET_0_73261, HIEFFPLA_NET_0_73262, 
        HIEFFPLA_NET_0_73263, HIEFFPLA_NET_0_73264, 
        HIEFFPLA_NET_0_73265, HIEFFPLA_NET_0_73266, 
        HIEFFPLA_NET_0_73267, HIEFFPLA_NET_0_73268, 
        HIEFFPLA_NET_0_73269, HIEFFPLA_NET_0_73270, 
        HIEFFPLA_NET_0_73271, HIEFFPLA_NET_0_73272, 
        HIEFFPLA_NET_0_73273, HIEFFPLA_NET_0_73274, 
        HIEFFPLA_NET_0_73275, HIEFFPLA_NET_0_73276, 
        HIEFFPLA_NET_0_73277, HIEFFPLA_NET_0_73278, 
        HIEFFPLA_NET_0_73279, HIEFFPLA_NET_0_73280, 
        HIEFFPLA_NET_0_73281, HIEFFPLA_NET_0_73282, 
        HIEFFPLA_NET_0_73283, HIEFFPLA_NET_0_73284, 
        HIEFFPLA_NET_0_73285, HIEFFPLA_NET_0_73286, 
        HIEFFPLA_NET_0_73287, HIEFFPLA_NET_0_73288, 
        HIEFFPLA_NET_0_73289, HIEFFPLA_NET_0_73290, 
        HIEFFPLA_NET_0_73291, HIEFFPLA_NET_0_73292, 
        HIEFFPLA_NET_0_73293, HIEFFPLA_NET_0_73294, 
        HIEFFPLA_NET_0_73295, HIEFFPLA_NET_0_73296, 
        HIEFFPLA_NET_0_73297, HIEFFPLA_NET_0_73298, 
        HIEFFPLA_NET_0_73299, HIEFFPLA_NET_0_73300, 
        HIEFFPLA_NET_0_73301, HIEFFPLA_NET_0_73302, 
        HIEFFPLA_NET_0_73303, HIEFFPLA_NET_0_73304, 
        HIEFFPLA_NET_0_73305, HIEFFPLA_NET_0_73306, 
        HIEFFPLA_NET_0_73307, HIEFFPLA_NET_0_73308, 
        HIEFFPLA_NET_0_73309, HIEFFPLA_NET_0_73310, 
        HIEFFPLA_NET_0_73311, HIEFFPLA_NET_0_73312, 
        HIEFFPLA_NET_0_73313, HIEFFPLA_NET_0_73314, 
        HIEFFPLA_NET_0_73315, HIEFFPLA_NET_0_73316, 
        HIEFFPLA_NET_0_73317, HIEFFPLA_NET_0_73318, 
        HIEFFPLA_NET_0_73319, HIEFFPLA_NET_0_73320, 
        HIEFFPLA_NET_0_73321, HIEFFPLA_NET_0_73322, 
        HIEFFPLA_NET_0_73323, HIEFFPLA_NET_0_73324, 
        HIEFFPLA_NET_0_73325, HIEFFPLA_NET_0_73326, 
        HIEFFPLA_NET_0_73327, HIEFFPLA_NET_0_73328, 
        HIEFFPLA_NET_0_73329, HIEFFPLA_NET_0_73330, 
        HIEFFPLA_NET_0_73331, HIEFFPLA_NET_0_73332, 
        HIEFFPLA_NET_0_73333, HIEFFPLA_NET_0_73334, 
        HIEFFPLA_NET_0_73335, HIEFFPLA_NET_0_73336, 
        HIEFFPLA_NET_0_73337, HIEFFPLA_NET_0_73338, 
        HIEFFPLA_NET_0_73339, HIEFFPLA_NET_0_73340, 
        HIEFFPLA_NET_0_73341, HIEFFPLA_NET_0_73342, 
        HIEFFPLA_NET_0_73343, HIEFFPLA_NET_0_73344, 
        HIEFFPLA_NET_0_73345, HIEFFPLA_NET_0_73346, 
        HIEFFPLA_NET_0_73347, HIEFFPLA_NET_0_73348, 
        HIEFFPLA_NET_0_73349, HIEFFPLA_NET_0_73350, 
        HIEFFPLA_NET_0_73351, HIEFFPLA_NET_0_73352, 
        HIEFFPLA_NET_0_73353, HIEFFPLA_NET_0_73354, 
        HIEFFPLA_NET_0_73355, HIEFFPLA_NET_0_73356, 
        HIEFFPLA_NET_0_73357, HIEFFPLA_NET_0_73358, 
        HIEFFPLA_NET_0_73359, HIEFFPLA_NET_0_73360, 
        HIEFFPLA_NET_0_73361, HIEFFPLA_NET_0_73362, 
        HIEFFPLA_NET_0_73363, HIEFFPLA_NET_0_73364, 
        HIEFFPLA_NET_0_73365, HIEFFPLA_NET_0_73366, 
        HIEFFPLA_NET_0_73367, HIEFFPLA_NET_0_73368, 
        HIEFFPLA_NET_0_73369, HIEFFPLA_NET_0_73370, 
        HIEFFPLA_NET_0_73371, HIEFFPLA_NET_0_73372, 
        HIEFFPLA_NET_0_73373, HIEFFPLA_NET_0_73374, 
        HIEFFPLA_NET_0_73375, HIEFFPLA_NET_0_73376, 
        HIEFFPLA_NET_0_73377, HIEFFPLA_NET_0_73378, 
        HIEFFPLA_NET_0_73379, HIEFFPLA_NET_0_73380, 
        HIEFFPLA_NET_0_73381, HIEFFPLA_NET_0_73382, 
        HIEFFPLA_NET_0_73383, HIEFFPLA_NET_0_73384, 
        HIEFFPLA_NET_0_73385, HIEFFPLA_NET_0_73386, 
        HIEFFPLA_NET_0_73387, HIEFFPLA_NET_0_73388, 
        HIEFFPLA_NET_0_73389, HIEFFPLA_NET_0_73390, 
        HIEFFPLA_NET_0_73391, HIEFFPLA_NET_0_73392, 
        HIEFFPLA_NET_0_73393, HIEFFPLA_NET_0_73394, 
        HIEFFPLA_NET_0_73395, HIEFFPLA_NET_0_73396, 
        HIEFFPLA_NET_0_73397, HIEFFPLA_NET_0_73398, 
        HIEFFPLA_NET_0_73399, HIEFFPLA_NET_0_73400, 
        HIEFFPLA_NET_0_73401, HIEFFPLA_NET_0_73402, 
        HIEFFPLA_NET_0_73403, HIEFFPLA_NET_0_73404, 
        HIEFFPLA_NET_0_73405, HIEFFPLA_NET_0_73406, 
        HIEFFPLA_NET_0_73407, HIEFFPLA_NET_0_73408, 
        HIEFFPLA_NET_0_73409, HIEFFPLA_NET_0_73410, 
        HIEFFPLA_NET_0_73411, HIEFFPLA_NET_0_73412, 
        HIEFFPLA_NET_0_73413, HIEFFPLA_NET_0_73414, 
        HIEFFPLA_NET_0_73415, HIEFFPLA_NET_0_73416, 
        HIEFFPLA_NET_0_73417, HIEFFPLA_NET_0_73418, 
        HIEFFPLA_NET_0_73419, HIEFFPLA_NET_0_73420, 
        HIEFFPLA_NET_0_73421, HIEFFPLA_NET_0_73422, 
        HIEFFPLA_NET_0_73423, HIEFFPLA_NET_0_73424, 
        HIEFFPLA_NET_0_73425, HIEFFPLA_NET_0_73426, 
        HIEFFPLA_NET_0_73427, HIEFFPLA_NET_0_73428, 
        HIEFFPLA_NET_0_73429, HIEFFPLA_NET_0_73430, 
        HIEFFPLA_NET_0_73431, HIEFFPLA_NET_0_73432, 
        HIEFFPLA_NET_0_73433, HIEFFPLA_NET_0_73434, 
        HIEFFPLA_NET_0_73435, HIEFFPLA_NET_0_73436, 
        HIEFFPLA_NET_0_73437, HIEFFPLA_NET_0_73438, 
        HIEFFPLA_NET_0_73439, HIEFFPLA_NET_0_73440, 
        HIEFFPLA_NET_0_73441, HIEFFPLA_NET_0_73442, 
        HIEFFPLA_NET_0_73443, HIEFFPLA_NET_0_73444, 
        HIEFFPLA_NET_0_73445, HIEFFPLA_NET_0_73446, 
        HIEFFPLA_NET_0_73447, HIEFFPLA_NET_0_73448, 
        HIEFFPLA_NET_0_73449, HIEFFPLA_NET_0_73450, 
        HIEFFPLA_NET_0_73451, HIEFFPLA_NET_0_73452, 
        HIEFFPLA_NET_0_73453, HIEFFPLA_NET_0_73454, 
        HIEFFPLA_NET_0_73455, HIEFFPLA_NET_0_73456, 
        HIEFFPLA_NET_0_73457, HIEFFPLA_NET_0_73458, 
        HIEFFPLA_NET_0_73459, HIEFFPLA_NET_0_73460, 
        HIEFFPLA_NET_0_73461, HIEFFPLA_NET_0_73462, 
        HIEFFPLA_NET_0_73463, HIEFFPLA_NET_0_73464, 
        HIEFFPLA_NET_0_73465, HIEFFPLA_NET_0_73466, 
        HIEFFPLA_NET_0_73467, HIEFFPLA_NET_0_73468, 
        HIEFFPLA_NET_0_73469, HIEFFPLA_NET_0_73470, 
        HIEFFPLA_NET_0_73471, HIEFFPLA_NET_0_73472, 
        HIEFFPLA_NET_0_73473, HIEFFPLA_NET_0_73474, 
        HIEFFPLA_NET_0_73475, HIEFFPLA_NET_0_73476, 
        HIEFFPLA_NET_0_73477, HIEFFPLA_NET_0_73478, 
        HIEFFPLA_NET_0_73479, HIEFFPLA_NET_0_73480, 
        HIEFFPLA_NET_0_73481, HIEFFPLA_NET_0_73482, 
        HIEFFPLA_NET_0_73483, HIEFFPLA_NET_0_73484, 
        HIEFFPLA_NET_0_73485, HIEFFPLA_NET_0_73486, 
        HIEFFPLA_NET_0_73487, HIEFFPLA_NET_0_73488, 
        HIEFFPLA_NET_0_73489, HIEFFPLA_NET_0_73490, 
        HIEFFPLA_NET_0_73491, HIEFFPLA_NET_0_73492, 
        HIEFFPLA_NET_0_73493, HIEFFPLA_NET_0_73494, 
        HIEFFPLA_NET_0_73495, HIEFFPLA_NET_0_73496, 
        HIEFFPLA_NET_0_73497, HIEFFPLA_NET_0_73498, 
        HIEFFPLA_NET_0_73499, HIEFFPLA_NET_0_73500, 
        HIEFFPLA_NET_0_73501, HIEFFPLA_NET_0_73502, 
        HIEFFPLA_NET_0_73503, HIEFFPLA_NET_0_73504, 
        HIEFFPLA_NET_0_73505, HIEFFPLA_NET_0_73506, 
        HIEFFPLA_NET_0_73507, HIEFFPLA_NET_0_73508, 
        HIEFFPLA_NET_0_73509, HIEFFPLA_NET_0_73510, 
        HIEFFPLA_NET_0_73511, HIEFFPLA_NET_0_73512, 
        HIEFFPLA_NET_0_73513, HIEFFPLA_NET_0_73514, 
        HIEFFPLA_NET_0_73515, HIEFFPLA_NET_0_73516, 
        HIEFFPLA_NET_0_73517, HIEFFPLA_NET_0_73518, 
        HIEFFPLA_NET_0_73519, HIEFFPLA_NET_0_73520, 
        HIEFFPLA_NET_0_73521, HIEFFPLA_NET_0_73522, 
        HIEFFPLA_NET_0_73523, HIEFFPLA_NET_0_73524, 
        HIEFFPLA_NET_0_73525, HIEFFPLA_NET_0_73526, 
        HIEFFPLA_NET_0_73527, HIEFFPLA_NET_0_73528, 
        HIEFFPLA_NET_0_73529, HIEFFPLA_NET_0_73530, 
        HIEFFPLA_NET_0_73531, HIEFFPLA_NET_0_73532, 
        HIEFFPLA_NET_0_73533, HIEFFPLA_NET_0_73534, 
        HIEFFPLA_NET_0_73535, HIEFFPLA_NET_0_73536, 
        HIEFFPLA_NET_0_73537, HIEFFPLA_NET_0_73538, 
        HIEFFPLA_NET_0_73539, HIEFFPLA_NET_0_73540, 
        HIEFFPLA_NET_0_73541, HIEFFPLA_NET_0_73542, 
        HIEFFPLA_NET_0_73543, HIEFFPLA_NET_0_73544, 
        HIEFFPLA_NET_0_73545, HIEFFPLA_NET_0_73546, 
        HIEFFPLA_NET_0_73547, HIEFFPLA_NET_0_73548, 
        HIEFFPLA_NET_0_73549, HIEFFPLA_NET_0_73550, 
        HIEFFPLA_NET_0_73551, HIEFFPLA_NET_0_73552, 
        HIEFFPLA_NET_0_73553, HIEFFPLA_NET_0_73554, 
        HIEFFPLA_NET_0_73555, HIEFFPLA_NET_0_73556, 
        HIEFFPLA_NET_0_73557, HIEFFPLA_NET_0_73558, 
        HIEFFPLA_NET_0_73559, HIEFFPLA_NET_0_73560, 
        HIEFFPLA_NET_0_73561, HIEFFPLA_NET_0_73562, 
        HIEFFPLA_NET_0_73563, HIEFFPLA_NET_0_73564, 
        HIEFFPLA_NET_0_73565, HIEFFPLA_NET_0_73566, 
        HIEFFPLA_NET_0_73567, HIEFFPLA_NET_0_73568, 
        HIEFFPLA_NET_0_73569, HIEFFPLA_NET_0_73570, 
        HIEFFPLA_NET_0_73571, HIEFFPLA_NET_0_73572, 
        HIEFFPLA_NET_0_73573, HIEFFPLA_NET_0_73574, 
        HIEFFPLA_NET_0_73575, HIEFFPLA_NET_0_73576, 
        HIEFFPLA_NET_0_73577, HIEFFPLA_NET_0_73578, 
        HIEFFPLA_NET_0_73579, HIEFFPLA_NET_0_73580, 
        HIEFFPLA_NET_0_73581, HIEFFPLA_NET_0_73582, 
        HIEFFPLA_NET_0_73583, HIEFFPLA_NET_0_73584, 
        HIEFFPLA_NET_0_73585, HIEFFPLA_NET_0_73586, 
        HIEFFPLA_NET_0_73587, HIEFFPLA_NET_0_73588, 
        HIEFFPLA_NET_0_73589, HIEFFPLA_NET_0_73590, 
        HIEFFPLA_NET_0_73591, HIEFFPLA_NET_0_73592, 
        HIEFFPLA_NET_0_73593, HIEFFPLA_NET_0_73594, 
        HIEFFPLA_NET_0_73595, HIEFFPLA_NET_0_73596, 
        HIEFFPLA_NET_0_73597, HIEFFPLA_NET_0_73598, 
        HIEFFPLA_NET_0_73599, HIEFFPLA_NET_0_73600, 
        HIEFFPLA_NET_0_73601, HIEFFPLA_NET_0_73602, 
        HIEFFPLA_NET_0_73603, HIEFFPLA_NET_0_73604, 
        HIEFFPLA_NET_0_73605, HIEFFPLA_NET_0_73606, 
        HIEFFPLA_NET_0_73607, HIEFFPLA_NET_0_73608, 
        HIEFFPLA_NET_0_73609, HIEFFPLA_NET_0_73610, 
        HIEFFPLA_NET_0_73611, HIEFFPLA_NET_0_73612, 
        HIEFFPLA_NET_0_73613, HIEFFPLA_NET_0_73614, 
        HIEFFPLA_NET_0_73615, HIEFFPLA_NET_0_73616, 
        HIEFFPLA_NET_0_73617, HIEFFPLA_NET_0_73618, 
        HIEFFPLA_NET_0_73619, HIEFFPLA_NET_0_73620, 
        HIEFFPLA_NET_0_73621, HIEFFPLA_NET_0_73622, 
        HIEFFPLA_NET_0_73623, HIEFFPLA_NET_0_73624, 
        HIEFFPLA_NET_0_73625, HIEFFPLA_NET_0_73626, 
        HIEFFPLA_NET_0_73627, HIEFFPLA_NET_0_73628, 
        HIEFFPLA_NET_0_73629, HIEFFPLA_NET_0_73630, 
        HIEFFPLA_NET_0_73631, HIEFFPLA_NET_0_73632, 
        HIEFFPLA_NET_0_73633, HIEFFPLA_NET_0_73634, 
        HIEFFPLA_NET_0_73635, HIEFFPLA_NET_0_73636, 
        HIEFFPLA_NET_0_73637, HIEFFPLA_NET_0_73638, 
        HIEFFPLA_NET_0_73639, HIEFFPLA_NET_0_73640, 
        HIEFFPLA_NET_0_73641, HIEFFPLA_NET_0_73642, 
        HIEFFPLA_NET_0_73643, HIEFFPLA_NET_0_73644, 
        HIEFFPLA_NET_0_73645, HIEFFPLA_NET_0_73646, 
        HIEFFPLA_NET_0_73647, HIEFFPLA_NET_0_73648, 
        HIEFFPLA_NET_0_73649, HIEFFPLA_NET_0_73650, 
        HIEFFPLA_NET_0_73651, HIEFFPLA_NET_0_73652, 
        HIEFFPLA_NET_0_73653, HIEFFPLA_NET_0_73654, 
        HIEFFPLA_NET_0_73655, HIEFFPLA_NET_0_73656, 
        HIEFFPLA_NET_0_73657, HIEFFPLA_NET_0_73658, 
        HIEFFPLA_NET_0_73659, HIEFFPLA_NET_0_73660, 
        HIEFFPLA_NET_0_73661, HIEFFPLA_NET_0_73662, 
        HIEFFPLA_NET_0_73663, HIEFFPLA_NET_0_73664, 
        HIEFFPLA_NET_0_73665, HIEFFPLA_NET_0_73666, 
        HIEFFPLA_NET_0_73667, HIEFFPLA_NET_0_73668, 
        HIEFFPLA_NET_0_73669, HIEFFPLA_NET_0_73670, 
        HIEFFPLA_NET_0_73671, HIEFFPLA_NET_0_73672, 
        HIEFFPLA_NET_0_73673, HIEFFPLA_NET_0_73674, 
        HIEFFPLA_NET_0_73675, HIEFFPLA_NET_0_73676, 
        HIEFFPLA_NET_0_73677, HIEFFPLA_NET_0_73678, 
        HIEFFPLA_NET_0_73679, HIEFFPLA_NET_0_73680, 
        HIEFFPLA_NET_0_73681, HIEFFPLA_NET_0_73682, 
        HIEFFPLA_NET_0_73683, HIEFFPLA_NET_0_73684, 
        HIEFFPLA_NET_0_73685, HIEFFPLA_NET_0_73686, 
        HIEFFPLA_NET_0_73687, HIEFFPLA_NET_0_73688, 
        HIEFFPLA_NET_0_73689, HIEFFPLA_NET_0_73690, 
        HIEFFPLA_NET_0_73691, HIEFFPLA_NET_0_73692, 
        HIEFFPLA_NET_0_73693, HIEFFPLA_NET_0_73694, 
        HIEFFPLA_NET_0_73695, HIEFFPLA_NET_0_73696, 
        HIEFFPLA_NET_0_73697, HIEFFPLA_NET_0_73698, 
        HIEFFPLA_NET_0_73699, HIEFFPLA_NET_0_73700, 
        HIEFFPLA_NET_0_73701, HIEFFPLA_NET_0_73702, 
        HIEFFPLA_NET_0_73703, HIEFFPLA_NET_0_73704, 
        HIEFFPLA_NET_0_73705, HIEFFPLA_NET_0_73706, 
        HIEFFPLA_NET_0_73707, HIEFFPLA_NET_0_73708, 
        HIEFFPLA_NET_0_73709, HIEFFPLA_NET_0_73710, 
        HIEFFPLA_NET_0_73711, HIEFFPLA_NET_0_73712, 
        HIEFFPLA_NET_0_73713, HIEFFPLA_NET_0_73714, 
        HIEFFPLA_NET_0_73715, HIEFFPLA_NET_0_73716, 
        HIEFFPLA_NET_0_73717, HIEFFPLA_NET_0_73718, 
        HIEFFPLA_NET_0_73719, HIEFFPLA_NET_0_73720, 
        HIEFFPLA_NET_0_73721, HIEFFPLA_NET_0_73722, 
        HIEFFPLA_NET_0_73723, HIEFFPLA_NET_0_73724, 
        HIEFFPLA_NET_0_73725, HIEFFPLA_NET_0_73726, 
        HIEFFPLA_NET_0_73727, HIEFFPLA_NET_0_73728, 
        HIEFFPLA_NET_0_73729, HIEFFPLA_NET_0_73730, 
        HIEFFPLA_NET_0_73731, HIEFFPLA_NET_0_73732, 
        HIEFFPLA_NET_0_73733, HIEFFPLA_NET_0_73734, 
        HIEFFPLA_NET_0_73735, HIEFFPLA_NET_0_73736, 
        HIEFFPLA_NET_0_73737, HIEFFPLA_NET_0_73738, 
        HIEFFPLA_NET_0_73739, HIEFFPLA_NET_0_73740, 
        HIEFFPLA_NET_0_73741, HIEFFPLA_NET_0_73742, 
        HIEFFPLA_NET_0_73743, HIEFFPLA_NET_0_73744, 
        HIEFFPLA_NET_0_73745, HIEFFPLA_NET_0_73746, 
        HIEFFPLA_NET_0_73747, HIEFFPLA_NET_0_73748, 
        HIEFFPLA_NET_0_73749, HIEFFPLA_NET_0_73750, 
        HIEFFPLA_NET_0_73751, HIEFFPLA_NET_0_73752, 
        HIEFFPLA_NET_0_73753, HIEFFPLA_NET_0_73754, 
        HIEFFPLA_NET_0_73755, HIEFFPLA_NET_0_73756, 
        HIEFFPLA_NET_0_73757, HIEFFPLA_NET_0_73758, 
        HIEFFPLA_NET_0_73759, HIEFFPLA_NET_0_73760, 
        HIEFFPLA_NET_0_73761, HIEFFPLA_NET_0_73762, 
        HIEFFPLA_NET_0_73763, HIEFFPLA_NET_0_73764, 
        HIEFFPLA_NET_0_73765, HIEFFPLA_NET_0_73766, 
        HIEFFPLA_NET_0_73767, HIEFFPLA_NET_0_73768, 
        HIEFFPLA_NET_0_73769, HIEFFPLA_NET_0_73770, 
        HIEFFPLA_NET_0_73771, HIEFFPLA_NET_0_73772, 
        HIEFFPLA_NET_0_73773, HIEFFPLA_NET_0_73774, 
        HIEFFPLA_NET_0_73775, HIEFFPLA_NET_0_73776, 
        HIEFFPLA_NET_0_73777, HIEFFPLA_NET_0_73778, 
        HIEFFPLA_NET_0_73779, HIEFFPLA_NET_0_73780, 
        HIEFFPLA_NET_0_73781, HIEFFPLA_NET_0_73782, 
        HIEFFPLA_NET_0_73783, HIEFFPLA_NET_0_73784, 
        HIEFFPLA_NET_0_73785, HIEFFPLA_NET_0_73786, 
        HIEFFPLA_NET_0_73787, HIEFFPLA_NET_0_73788, 
        HIEFFPLA_NET_0_73789, HIEFFPLA_NET_0_73790, 
        HIEFFPLA_NET_0_73791, HIEFFPLA_NET_0_73792, 
        HIEFFPLA_NET_0_73793, HIEFFPLA_NET_0_73794, 
        HIEFFPLA_NET_0_73795, HIEFFPLA_NET_0_73796, 
        HIEFFPLA_NET_0_73797, HIEFFPLA_NET_0_73798, 
        HIEFFPLA_NET_0_73799, HIEFFPLA_NET_0_73800, 
        HIEFFPLA_NET_0_73801, HIEFFPLA_NET_0_73802, 
        HIEFFPLA_NET_0_73803, HIEFFPLA_NET_0_73804, 
        HIEFFPLA_NET_0_73805, HIEFFPLA_NET_0_73806, 
        HIEFFPLA_NET_0_73807, HIEFFPLA_NET_0_73808, 
        HIEFFPLA_NET_0_73809, HIEFFPLA_NET_0_73810, 
        HIEFFPLA_NET_0_73811, HIEFFPLA_NET_0_73812, 
        HIEFFPLA_NET_0_73813, HIEFFPLA_NET_0_73814, 
        HIEFFPLA_NET_0_73815, HIEFFPLA_NET_0_73816, 
        HIEFFPLA_NET_0_73817, HIEFFPLA_NET_0_73818, 
        HIEFFPLA_NET_0_73819, HIEFFPLA_NET_0_73820, 
        HIEFFPLA_NET_0_73821, HIEFFPLA_NET_0_73822, 
        HIEFFPLA_NET_0_73823, HIEFFPLA_NET_0_73824, 
        HIEFFPLA_NET_0_73825, HIEFFPLA_NET_0_73826, 
        HIEFFPLA_NET_0_73827, HIEFFPLA_NET_0_73828, 
        HIEFFPLA_NET_0_73829, HIEFFPLA_NET_0_73830, 
        HIEFFPLA_NET_0_73831, HIEFFPLA_NET_0_73832, 
        HIEFFPLA_NET_0_73833, HIEFFPLA_NET_0_73834, 
        HIEFFPLA_NET_0_73835, HIEFFPLA_NET_0_73836, 
        HIEFFPLA_NET_0_73837, HIEFFPLA_NET_0_73838, 
        HIEFFPLA_NET_0_73839, HIEFFPLA_NET_0_73840, 
        HIEFFPLA_NET_0_73841, HIEFFPLA_NET_0_73842, 
        HIEFFPLA_NET_0_73843, HIEFFPLA_NET_0_73844, 
        HIEFFPLA_NET_0_73845, HIEFFPLA_NET_0_73846, 
        HIEFFPLA_NET_0_73847, HIEFFPLA_NET_0_73848, 
        HIEFFPLA_NET_0_73849, HIEFFPLA_NET_0_73850, 
        HIEFFPLA_NET_0_73851, HIEFFPLA_NET_0_73852, 
        HIEFFPLA_NET_0_73853, HIEFFPLA_NET_0_73854, 
        HIEFFPLA_NET_0_73855, HIEFFPLA_NET_0_73856, 
        HIEFFPLA_NET_0_73857, HIEFFPLA_NET_0_73858, 
        HIEFFPLA_NET_0_73859, HIEFFPLA_NET_0_73860, 
        HIEFFPLA_NET_0_73861, HIEFFPLA_NET_0_73862, 
        HIEFFPLA_NET_0_73863, HIEFFPLA_NET_0_73864, 
        HIEFFPLA_NET_0_73865, HIEFFPLA_NET_0_73866, 
        HIEFFPLA_NET_0_73867, HIEFFPLA_NET_0_73868, 
        HIEFFPLA_NET_0_73869, HIEFFPLA_NET_0_73870, 
        HIEFFPLA_NET_0_73871, HIEFFPLA_NET_0_73872, 
        HIEFFPLA_NET_0_73873, HIEFFPLA_NET_0_73874, 
        HIEFFPLA_NET_0_73875, HIEFFPLA_NET_0_73876, 
        HIEFFPLA_NET_0_73877, HIEFFPLA_NET_0_73878, 
        HIEFFPLA_NET_0_73879, HIEFFPLA_NET_0_73880, 
        HIEFFPLA_NET_0_73881, HIEFFPLA_NET_0_73882, 
        HIEFFPLA_NET_0_73883, HIEFFPLA_NET_0_73884, 
        HIEFFPLA_NET_0_73885, HIEFFPLA_NET_0_73886, 
        HIEFFPLA_NET_0_73887, HIEFFPLA_NET_0_73888, 
        HIEFFPLA_NET_0_73889, HIEFFPLA_NET_0_73890, 
        HIEFFPLA_NET_0_73891, HIEFFPLA_NET_0_73892, 
        HIEFFPLA_NET_0_73893, HIEFFPLA_NET_0_73894, 
        HIEFFPLA_NET_0_73895, HIEFFPLA_NET_0_73896, 
        HIEFFPLA_NET_0_73897, HIEFFPLA_NET_0_73898, 
        HIEFFPLA_NET_0_73899, HIEFFPLA_NET_0_73900, 
        HIEFFPLA_NET_0_73901, HIEFFPLA_NET_0_73902, 
        HIEFFPLA_NET_0_73903, HIEFFPLA_NET_0_73904, 
        HIEFFPLA_NET_0_73905, HIEFFPLA_NET_0_73906, 
        HIEFFPLA_NET_0_73907, HIEFFPLA_NET_0_73908, 
        HIEFFPLA_NET_0_73909, HIEFFPLA_NET_0_73910, 
        HIEFFPLA_NET_0_73911, HIEFFPLA_NET_0_73912, 
        HIEFFPLA_NET_0_73913, HIEFFPLA_NET_0_73914, 
        HIEFFPLA_NET_0_73915, HIEFFPLA_NET_0_73916, 
        HIEFFPLA_NET_0_73917, HIEFFPLA_NET_0_73918, 
        HIEFFPLA_NET_0_73919, HIEFFPLA_NET_0_73920, 
        HIEFFPLA_NET_0_73921, HIEFFPLA_NET_0_73922, 
        HIEFFPLA_NET_0_73923, HIEFFPLA_NET_0_73924, 
        HIEFFPLA_NET_0_73925, HIEFFPLA_NET_0_73926, 
        HIEFFPLA_NET_0_73927, HIEFFPLA_NET_0_73928, 
        HIEFFPLA_NET_0_73929, HIEFFPLA_NET_0_73930, 
        HIEFFPLA_NET_0_73931, HIEFFPLA_NET_0_73932, 
        HIEFFPLA_NET_0_73933, HIEFFPLA_NET_0_73934, 
        HIEFFPLA_NET_0_73935, HIEFFPLA_NET_0_73936, 
        HIEFFPLA_NET_0_73937, HIEFFPLA_NET_0_73938, 
        HIEFFPLA_NET_0_73939, HIEFFPLA_NET_0_73940, 
        HIEFFPLA_NET_0_73941, HIEFFPLA_NET_0_73942, 
        HIEFFPLA_NET_0_73943, HIEFFPLA_NET_0_73944, 
        HIEFFPLA_NET_0_73945, HIEFFPLA_NET_0_73946, 
        HIEFFPLA_NET_0_73947, HIEFFPLA_NET_0_73948, 
        HIEFFPLA_NET_0_73949, HIEFFPLA_NET_0_73950, 
        HIEFFPLA_NET_0_73951, HIEFFPLA_NET_0_73952, 
        HIEFFPLA_NET_0_73953, HIEFFPLA_NET_0_73954, 
        HIEFFPLA_NET_0_73955, HIEFFPLA_NET_0_73956, 
        HIEFFPLA_NET_0_73957, HIEFFPLA_NET_0_73958, 
        HIEFFPLA_NET_0_73959, HIEFFPLA_NET_0_73960, 
        HIEFFPLA_NET_0_73961, HIEFFPLA_NET_0_73962, 
        HIEFFPLA_NET_0_73963, HIEFFPLA_NET_0_73964, 
        HIEFFPLA_NET_0_73965, HIEFFPLA_NET_0_73966, 
        HIEFFPLA_NET_0_73967, HIEFFPLA_NET_0_73968, 
        HIEFFPLA_NET_0_73969, HIEFFPLA_NET_0_73970, 
        HIEFFPLA_NET_0_73971, HIEFFPLA_NET_0_73972, 
        HIEFFPLA_NET_0_73973, HIEFFPLA_NET_0_73974, 
        HIEFFPLA_NET_0_73975, HIEFFPLA_NET_0_73976, 
        HIEFFPLA_NET_0_73977, HIEFFPLA_NET_0_73978, 
        HIEFFPLA_NET_0_73979, HIEFFPLA_NET_0_73980, 
        HIEFFPLA_NET_0_73981, HIEFFPLA_NET_0_73982, 
        HIEFFPLA_NET_0_73983, HIEFFPLA_NET_0_73984, 
        HIEFFPLA_NET_0_73985, HIEFFPLA_NET_0_73986, 
        HIEFFPLA_NET_0_73987, HIEFFPLA_NET_0_73988, 
        HIEFFPLA_NET_0_73989, HIEFFPLA_NET_0_73990, 
        HIEFFPLA_NET_0_73991, HIEFFPLA_NET_0_73992, 
        HIEFFPLA_NET_0_73993, HIEFFPLA_NET_0_73994, 
        HIEFFPLA_NET_0_73995, HIEFFPLA_NET_0_73996, 
        HIEFFPLA_NET_0_73997, HIEFFPLA_NET_0_73998, 
        HIEFFPLA_NET_0_73999, HIEFFPLA_NET_0_74000, 
        HIEFFPLA_NET_0_74001, HIEFFPLA_NET_0_74002, 
        HIEFFPLA_NET_0_74003, HIEFFPLA_NET_0_74004, 
        HIEFFPLA_NET_0_74005, HIEFFPLA_NET_0_74006, 
        HIEFFPLA_NET_0_74007, HIEFFPLA_NET_0_74008, 
        HIEFFPLA_NET_0_74009, HIEFFPLA_NET_0_74010, 
        HIEFFPLA_NET_0_74011, HIEFFPLA_NET_0_74012, 
        HIEFFPLA_NET_0_74013, HIEFFPLA_NET_0_74014, 
        HIEFFPLA_NET_0_74015, HIEFFPLA_NET_0_74016, 
        HIEFFPLA_NET_0_74017, HIEFFPLA_NET_0_74018, 
        HIEFFPLA_NET_0_74019, HIEFFPLA_NET_0_74020, 
        HIEFFPLA_NET_0_74021, HIEFFPLA_NET_0_74022, 
        HIEFFPLA_NET_0_74023, HIEFFPLA_NET_0_74024, 
        HIEFFPLA_NET_0_74025, HIEFFPLA_NET_0_74026, 
        HIEFFPLA_NET_0_74027, HIEFFPLA_NET_0_74028, 
        HIEFFPLA_NET_0_74029, HIEFFPLA_NET_0_74030, 
        HIEFFPLA_NET_0_74031, HIEFFPLA_NET_0_74032, 
        HIEFFPLA_NET_0_74033, HIEFFPLA_NET_0_74034, 
        HIEFFPLA_NET_0_74035, HIEFFPLA_NET_0_74036, 
        HIEFFPLA_NET_0_74037, HIEFFPLA_NET_0_74038, 
        HIEFFPLA_NET_0_74039, HIEFFPLA_NET_0_74040, 
        HIEFFPLA_NET_0_74041, HIEFFPLA_NET_0_74042, 
        HIEFFPLA_NET_0_74043, HIEFFPLA_NET_0_74044, 
        HIEFFPLA_NET_0_74045, HIEFFPLA_NET_0_74046, 
        HIEFFPLA_NET_0_74047, HIEFFPLA_NET_0_74048, 
        HIEFFPLA_NET_0_74049, HIEFFPLA_NET_0_74050, 
        HIEFFPLA_NET_0_74051, HIEFFPLA_NET_0_74052, 
        HIEFFPLA_NET_0_74053, HIEFFPLA_NET_0_74054, 
        HIEFFPLA_NET_0_74055, HIEFFPLA_NET_0_74056, 
        HIEFFPLA_NET_0_74057, HIEFFPLA_NET_0_74058, 
        HIEFFPLA_NET_0_74059, HIEFFPLA_NET_0_74060, 
        HIEFFPLA_NET_0_74061, HIEFFPLA_NET_0_74062, 
        HIEFFPLA_NET_0_74063, HIEFFPLA_NET_0_74064, 
        HIEFFPLA_NET_0_74065, HIEFFPLA_NET_0_74066, 
        HIEFFPLA_NET_0_74067, HIEFFPLA_NET_0_74068, 
        HIEFFPLA_NET_0_74069, HIEFFPLA_NET_0_74070, 
        HIEFFPLA_NET_0_74071, HIEFFPLA_NET_0_74072, 
        HIEFFPLA_NET_0_74073, HIEFFPLA_NET_0_74074, 
        HIEFFPLA_NET_0_74075, HIEFFPLA_NET_0_74076, 
        HIEFFPLA_NET_0_74077, HIEFFPLA_NET_0_74078, 
        HIEFFPLA_NET_0_74079, HIEFFPLA_NET_0_74080, 
        HIEFFPLA_NET_0_74081, HIEFFPLA_NET_0_74082, 
        HIEFFPLA_NET_0_74083, HIEFFPLA_NET_0_74084, 
        HIEFFPLA_NET_0_74085, HIEFFPLA_NET_0_74086, 
        HIEFFPLA_NET_0_74087, HIEFFPLA_NET_0_74088, 
        HIEFFPLA_NET_0_74089, HIEFFPLA_NET_0_74090, 
        HIEFFPLA_NET_0_74091, HIEFFPLA_NET_0_74092, 
        HIEFFPLA_NET_0_74093, HIEFFPLA_NET_0_74094, 
        HIEFFPLA_NET_0_74095, HIEFFPLA_NET_0_74096, 
        HIEFFPLA_NET_0_74097, HIEFFPLA_NET_0_74098, 
        HIEFFPLA_NET_0_74099, HIEFFPLA_NET_0_74100, 
        HIEFFPLA_NET_0_74101, HIEFFPLA_NET_0_74102, 
        HIEFFPLA_NET_0_74103, HIEFFPLA_NET_0_74104, 
        HIEFFPLA_NET_0_74105, HIEFFPLA_NET_0_74106, 
        HIEFFPLA_NET_0_74107, HIEFFPLA_NET_0_74108, 
        HIEFFPLA_NET_0_74109, HIEFFPLA_NET_0_74110, 
        HIEFFPLA_NET_0_74111, HIEFFPLA_NET_0_74112, 
        HIEFFPLA_NET_0_74113, HIEFFPLA_NET_0_74114, 
        HIEFFPLA_NET_0_74115, HIEFFPLA_NET_0_74116, 
        HIEFFPLA_NET_0_74117, HIEFFPLA_NET_0_74118, 
        HIEFFPLA_NET_0_74119, HIEFFPLA_NET_0_74120, 
        HIEFFPLA_NET_0_74121, HIEFFPLA_NET_0_74122, 
        HIEFFPLA_NET_0_74123, HIEFFPLA_NET_0_74124, 
        HIEFFPLA_NET_0_74125, HIEFFPLA_NET_0_74126, 
        HIEFFPLA_NET_0_74127, HIEFFPLA_NET_0_74128, 
        HIEFFPLA_NET_0_74129, HIEFFPLA_NET_0_74130, 
        HIEFFPLA_NET_0_74131, HIEFFPLA_NET_0_74132, 
        HIEFFPLA_NET_0_74133, HIEFFPLA_NET_0_74134, 
        HIEFFPLA_NET_0_74135, HIEFFPLA_NET_0_74136, 
        HIEFFPLA_NET_0_74137, HIEFFPLA_NET_0_74138, 
        HIEFFPLA_NET_0_74139, HIEFFPLA_NET_0_74140, 
        HIEFFPLA_NET_0_74141, HIEFFPLA_NET_0_74142, 
        HIEFFPLA_NET_0_74143, HIEFFPLA_NET_0_74144, 
        HIEFFPLA_NET_0_74145, HIEFFPLA_NET_0_74146, 
        HIEFFPLA_NET_0_74147, HIEFFPLA_NET_0_74148, 
        HIEFFPLA_NET_0_74149, HIEFFPLA_NET_0_74150, 
        HIEFFPLA_NET_0_74151, HIEFFPLA_NET_0_74152, 
        HIEFFPLA_NET_0_74153, HIEFFPLA_NET_0_74154, 
        HIEFFPLA_NET_0_74155, HIEFFPLA_NET_0_74156, 
        HIEFFPLA_NET_0_74157, HIEFFPLA_NET_0_74158, 
        HIEFFPLA_NET_0_74159, HIEFFPLA_NET_0_74160, 
        HIEFFPLA_NET_0_74161, HIEFFPLA_NET_0_74162, 
        HIEFFPLA_NET_0_74163, HIEFFPLA_NET_0_74164, 
        HIEFFPLA_NET_0_74165, HIEFFPLA_NET_0_74166, 
        HIEFFPLA_NET_0_74167, HIEFFPLA_NET_0_74168, 
        HIEFFPLA_NET_0_74169, HIEFFPLA_NET_0_74170, 
        HIEFFPLA_NET_0_74171, HIEFFPLA_NET_0_74172, 
        HIEFFPLA_NET_0_74173, HIEFFPLA_NET_0_74174, 
        HIEFFPLA_NET_0_74175, HIEFFPLA_NET_0_74176, 
        HIEFFPLA_NET_0_74177, HIEFFPLA_NET_0_74178, 
        HIEFFPLA_NET_0_74179, HIEFFPLA_NET_0_74180, 
        HIEFFPLA_NET_0_74181, HIEFFPLA_NET_0_74182, 
        HIEFFPLA_NET_0_74183, HIEFFPLA_NET_0_74184, 
        HIEFFPLA_NET_0_74185, HIEFFPLA_NET_0_74186, 
        HIEFFPLA_NET_0_74187, HIEFFPLA_NET_0_74188, 
        HIEFFPLA_NET_0_74189, HIEFFPLA_NET_0_74190, 
        HIEFFPLA_NET_0_74191, HIEFFPLA_NET_0_74192, 
        HIEFFPLA_NET_0_74193, HIEFFPLA_NET_0_74194, 
        HIEFFPLA_NET_0_74195, HIEFFPLA_NET_0_74196, 
        HIEFFPLA_NET_0_74197, HIEFFPLA_NET_0_74198, 
        HIEFFPLA_NET_0_74199, HIEFFPLA_NET_0_74200, 
        HIEFFPLA_NET_0_74201, HIEFFPLA_NET_0_74202, 
        HIEFFPLA_NET_0_74203, HIEFFPLA_NET_0_74204, 
        HIEFFPLA_NET_0_74205, HIEFFPLA_NET_0_74206, 
        HIEFFPLA_NET_0_74207, HIEFFPLA_NET_0_74208, 
        HIEFFPLA_NET_0_74209, HIEFFPLA_NET_0_74210, 
        HIEFFPLA_NET_0_74211, HIEFFPLA_NET_0_74212, 
        HIEFFPLA_NET_0_74213, HIEFFPLA_NET_0_74214, 
        HIEFFPLA_NET_0_74215, HIEFFPLA_NET_0_74216, 
        HIEFFPLA_NET_0_74217, HIEFFPLA_NET_0_74218, 
        HIEFFPLA_NET_0_74219, HIEFFPLA_NET_0_74220, 
        HIEFFPLA_NET_0_74221, HIEFFPLA_NET_0_74222, 
        HIEFFPLA_NET_0_74223, HIEFFPLA_NET_0_74224, 
        HIEFFPLA_NET_0_74225, HIEFFPLA_NET_0_74226, 
        HIEFFPLA_NET_0_74227, HIEFFPLA_NET_0_74228, 
        HIEFFPLA_NET_0_74229, HIEFFPLA_NET_0_74230, 
        HIEFFPLA_NET_0_74231, HIEFFPLA_NET_0_74232, 
        HIEFFPLA_NET_0_74233, HIEFFPLA_NET_0_74234, 
        HIEFFPLA_NET_0_74235, HIEFFPLA_NET_0_74236, 
        HIEFFPLA_NET_0_74237, HIEFFPLA_NET_0_74238, 
        HIEFFPLA_NET_0_74239, HIEFFPLA_NET_0_74240, 
        HIEFFPLA_NET_0_74241, HIEFFPLA_NET_0_74242, 
        HIEFFPLA_NET_0_74243, HIEFFPLA_NET_0_74244, 
        HIEFFPLA_NET_0_74245, HIEFFPLA_NET_0_74246, 
        HIEFFPLA_NET_0_74247, HIEFFPLA_NET_0_74248, 
        HIEFFPLA_NET_0_74249, HIEFFPLA_NET_0_74250, 
        HIEFFPLA_NET_0_74251, HIEFFPLA_NET_0_74252, 
        HIEFFPLA_NET_0_74253, HIEFFPLA_NET_0_74254, 
        HIEFFPLA_NET_0_74255, HIEFFPLA_NET_0_74256, 
        HIEFFPLA_NET_0_74257, HIEFFPLA_NET_0_74258, 
        HIEFFPLA_NET_0_74259, HIEFFPLA_NET_0_74260, 
        HIEFFPLA_NET_0_74261, HIEFFPLA_NET_0_74262, 
        HIEFFPLA_NET_0_74263, HIEFFPLA_NET_0_74264, 
        HIEFFPLA_NET_0_74265, HIEFFPLA_NET_0_74266, 
        HIEFFPLA_NET_0_74267, HIEFFPLA_NET_0_74268, 
        HIEFFPLA_NET_0_74269, HIEFFPLA_NET_0_74270, 
        HIEFFPLA_NET_0_74271, HIEFFPLA_NET_0_74272, 
        HIEFFPLA_NET_0_74273, HIEFFPLA_NET_0_74274, 
        HIEFFPLA_NET_0_74275, HIEFFPLA_NET_0_74276, 
        HIEFFPLA_NET_0_74277, HIEFFPLA_NET_0_74278, 
        HIEFFPLA_NET_0_74279, HIEFFPLA_NET_0_74280, 
        HIEFFPLA_NET_0_74281, HIEFFPLA_NET_0_74282, 
        HIEFFPLA_NET_0_74283, HIEFFPLA_NET_0_74284, 
        HIEFFPLA_NET_0_74285, HIEFFPLA_NET_0_74286, 
        HIEFFPLA_NET_0_74287, HIEFFPLA_NET_0_74288, 
        HIEFFPLA_NET_0_74289, HIEFFPLA_NET_0_74290, 
        HIEFFPLA_NET_0_74291, HIEFFPLA_NET_0_74292, 
        HIEFFPLA_NET_0_74293, HIEFFPLA_NET_0_74294, 
        HIEFFPLA_NET_0_74295, HIEFFPLA_NET_0_74296, 
        HIEFFPLA_NET_0_74297, HIEFFPLA_NET_0_74298, 
        HIEFFPLA_NET_0_74299, HIEFFPLA_NET_0_74300, 
        HIEFFPLA_NET_0_74301, HIEFFPLA_NET_0_74302, 
        HIEFFPLA_NET_0_74303, HIEFFPLA_NET_0_74304, 
        HIEFFPLA_NET_0_74305, HIEFFPLA_NET_0_74306, 
        HIEFFPLA_NET_0_74307, HIEFFPLA_NET_0_74308, 
        HIEFFPLA_NET_0_74309, HIEFFPLA_NET_0_74310, 
        HIEFFPLA_NET_0_74311, HIEFFPLA_NET_0_74312, 
        HIEFFPLA_NET_0_74313, HIEFFPLA_NET_0_74314, 
        HIEFFPLA_NET_0_74315, HIEFFPLA_NET_0_74316, 
        HIEFFPLA_NET_0_74317, HIEFFPLA_NET_0_74318, 
        HIEFFPLA_NET_0_74319, HIEFFPLA_NET_0_74320, 
        HIEFFPLA_NET_0_74321, HIEFFPLA_NET_0_74322, 
        HIEFFPLA_NET_0_74323, HIEFFPLA_NET_0_74324, 
        HIEFFPLA_NET_0_74325, HIEFFPLA_NET_0_74326, 
        HIEFFPLA_NET_0_74327, HIEFFPLA_NET_0_74328, 
        HIEFFPLA_NET_0_74329, HIEFFPLA_NET_0_74330, 
        HIEFFPLA_NET_0_74331, HIEFFPLA_NET_0_74332, 
        HIEFFPLA_NET_0_74333, HIEFFPLA_NET_0_74334, 
        HIEFFPLA_NET_0_74335, HIEFFPLA_NET_0_74336, 
        HIEFFPLA_NET_0_74337, HIEFFPLA_NET_0_74338, 
        HIEFFPLA_NET_0_74339, HIEFFPLA_NET_0_74340, 
        HIEFFPLA_NET_0_74341, HIEFFPLA_NET_0_74342, 
        HIEFFPLA_NET_0_74343, HIEFFPLA_NET_0_74344, 
        HIEFFPLA_NET_0_74345, HIEFFPLA_NET_0_74346, 
        HIEFFPLA_NET_0_74347, HIEFFPLA_NET_0_74348, 
        HIEFFPLA_NET_0_74349, HIEFFPLA_NET_0_74350, 
        HIEFFPLA_NET_0_74351, HIEFFPLA_NET_0_74352, 
        HIEFFPLA_NET_0_74353, HIEFFPLA_NET_0_74354, 
        HIEFFPLA_NET_0_74355, HIEFFPLA_NET_0_74356, 
        HIEFFPLA_NET_0_74357, HIEFFPLA_NET_0_74358, 
        HIEFFPLA_NET_0_74359, HIEFFPLA_NET_0_74360, 
        HIEFFPLA_NET_0_74361, HIEFFPLA_NET_0_74362, 
        HIEFFPLA_NET_0_74363, HIEFFPLA_NET_0_74364, 
        HIEFFPLA_NET_0_74365, HIEFFPLA_NET_0_74366, 
        HIEFFPLA_NET_0_74367, HIEFFPLA_NET_0_74368, 
        HIEFFPLA_NET_0_74369, HIEFFPLA_NET_0_74370, 
        HIEFFPLA_NET_0_74371, HIEFFPLA_NET_0_74372, 
        HIEFFPLA_NET_0_74373, HIEFFPLA_NET_0_74374, 
        HIEFFPLA_NET_0_74375, HIEFFPLA_NET_0_74376, 
        HIEFFPLA_NET_0_74377, HIEFFPLA_NET_0_74378, 
        HIEFFPLA_NET_0_74379, HIEFFPLA_NET_0_74380, 
        HIEFFPLA_NET_0_74381, HIEFFPLA_NET_0_74382, 
        HIEFFPLA_NET_0_74383, HIEFFPLA_NET_0_74384, 
        HIEFFPLA_NET_0_74385, HIEFFPLA_NET_0_74386, 
        HIEFFPLA_NET_0_74387, HIEFFPLA_NET_0_74388, 
        HIEFFPLA_NET_0_74389, HIEFFPLA_NET_0_74390, 
        HIEFFPLA_NET_0_74391, HIEFFPLA_NET_0_74392, 
        HIEFFPLA_NET_0_74393, HIEFFPLA_NET_0_74394, 
        HIEFFPLA_NET_0_74395, HIEFFPLA_NET_0_74396, 
        HIEFFPLA_NET_0_74397, HIEFFPLA_NET_0_74398, 
        HIEFFPLA_NET_0_74399, HIEFFPLA_NET_0_74400, 
        HIEFFPLA_NET_0_74401, HIEFFPLA_NET_0_74402, 
        HIEFFPLA_NET_0_74403, HIEFFPLA_NET_0_74404, 
        HIEFFPLA_NET_0_74405, HIEFFPLA_NET_0_74406, 
        HIEFFPLA_NET_0_74407, HIEFFPLA_NET_0_74408, 
        HIEFFPLA_NET_0_74409, HIEFFPLA_NET_0_74410, 
        HIEFFPLA_NET_0_74411, HIEFFPLA_NET_0_74412, 
        HIEFFPLA_NET_0_74413, HIEFFPLA_NET_0_74414, 
        HIEFFPLA_NET_0_74415, HIEFFPLA_NET_0_74416, 
        HIEFFPLA_NET_0_74417, HIEFFPLA_NET_0_74418, 
        HIEFFPLA_NET_0_74419, HIEFFPLA_NET_0_74420, 
        HIEFFPLA_NET_0_74421, HIEFFPLA_NET_0_74422, 
        HIEFFPLA_NET_0_74423, HIEFFPLA_NET_0_74424, 
        HIEFFPLA_NET_0_74425, HIEFFPLA_NET_0_74426, 
        HIEFFPLA_NET_0_74427, HIEFFPLA_NET_0_74428, 
        HIEFFPLA_NET_0_74429, HIEFFPLA_NET_0_74430, 
        HIEFFPLA_NET_0_74431, HIEFFPLA_NET_0_74432, 
        HIEFFPLA_NET_0_74433, HIEFFPLA_NET_0_74434, 
        HIEFFPLA_NET_0_74435, HIEFFPLA_NET_0_74436, 
        HIEFFPLA_NET_0_74437, HIEFFPLA_NET_0_74438, 
        HIEFFPLA_NET_0_74439, HIEFFPLA_NET_0_74440, 
        HIEFFPLA_NET_0_74441, HIEFFPLA_NET_0_74442, 
        HIEFFPLA_NET_0_74443, HIEFFPLA_NET_0_74444, 
        HIEFFPLA_NET_0_74445, HIEFFPLA_NET_0_74446, 
        HIEFFPLA_NET_0_74447, HIEFFPLA_NET_0_74448, 
        HIEFFPLA_NET_0_74449, HIEFFPLA_NET_0_74450, 
        HIEFFPLA_NET_0_74451, HIEFFPLA_NET_0_74452, 
        HIEFFPLA_NET_0_74453, HIEFFPLA_NET_0_74454, 
        HIEFFPLA_NET_0_74455, HIEFFPLA_NET_0_74456, 
        HIEFFPLA_NET_0_74457, HIEFFPLA_NET_0_74458, 
        HIEFFPLA_NET_0_74459, HIEFFPLA_NET_0_74460, 
        HIEFFPLA_NET_0_74461, HIEFFPLA_NET_0_74462, 
        HIEFFPLA_NET_0_74463, HIEFFPLA_NET_0_74464, 
        HIEFFPLA_NET_0_74465, HIEFFPLA_NET_0_74466, 
        HIEFFPLA_NET_0_74467, HIEFFPLA_NET_0_74468, 
        HIEFFPLA_NET_0_74469, HIEFFPLA_NET_0_74470, 
        HIEFFPLA_NET_0_74471, HIEFFPLA_NET_0_74472, 
        HIEFFPLA_NET_0_74473, HIEFFPLA_NET_0_74474, 
        HIEFFPLA_NET_0_74475, HIEFFPLA_NET_0_74476, 
        HIEFFPLA_NET_0_74477, HIEFFPLA_NET_0_74478, 
        HIEFFPLA_NET_0_74479, HIEFFPLA_NET_0_74480, 
        HIEFFPLA_NET_0_74481, HIEFFPLA_NET_0_74482, 
        HIEFFPLA_NET_0_74483, HIEFFPLA_NET_0_74484, 
        HIEFFPLA_NET_0_74485, HIEFFPLA_NET_0_74486, 
        HIEFFPLA_NET_0_74487, HIEFFPLA_NET_0_74488, 
        HIEFFPLA_NET_0_74489, HIEFFPLA_NET_0_74490, 
        HIEFFPLA_NET_0_74491, HIEFFPLA_NET_0_74492, 
        HIEFFPLA_NET_0_74493, HIEFFPLA_NET_0_74494, 
        HIEFFPLA_NET_0_74495, HIEFFPLA_NET_0_74496, 
        HIEFFPLA_NET_0_74497, HIEFFPLA_NET_0_74498, 
        HIEFFPLA_NET_0_74499, HIEFFPLA_NET_0_74500, 
        HIEFFPLA_NET_0_74501, HIEFFPLA_NET_0_74502, 
        HIEFFPLA_NET_0_74503, HIEFFPLA_NET_0_74504, 
        HIEFFPLA_NET_0_74505, HIEFFPLA_NET_0_74506, 
        HIEFFPLA_NET_0_74507, HIEFFPLA_NET_0_74508, 
        HIEFFPLA_NET_0_74509, HIEFFPLA_NET_0_74510, 
        HIEFFPLA_NET_0_74511, HIEFFPLA_NET_0_74512, 
        HIEFFPLA_NET_0_74513, HIEFFPLA_NET_0_74514, 
        HIEFFPLA_NET_0_74515, HIEFFPLA_NET_0_74516, 
        HIEFFPLA_NET_0_74517, HIEFFPLA_NET_0_74518, 
        HIEFFPLA_NET_0_74519, HIEFFPLA_NET_0_74520, 
        HIEFFPLA_NET_0_74521, HIEFFPLA_NET_0_74522, 
        HIEFFPLA_NET_0_74523, HIEFFPLA_NET_0_74524, 
        HIEFFPLA_NET_0_74525, HIEFFPLA_NET_0_74526, 
        HIEFFPLA_NET_0_74527, HIEFFPLA_NET_0_74528, 
        HIEFFPLA_NET_0_74529, HIEFFPLA_NET_0_74530, 
        HIEFFPLA_NET_0_74531, HIEFFPLA_NET_0_74532, 
        HIEFFPLA_NET_0_74533, HIEFFPLA_NET_0_74534, 
        HIEFFPLA_NET_0_74535, HIEFFPLA_NET_0_74536, 
        HIEFFPLA_NET_0_74537, HIEFFPLA_NET_0_74538, 
        HIEFFPLA_NET_0_74539, HIEFFPLA_NET_0_74540, 
        HIEFFPLA_NET_0_74541, HIEFFPLA_NET_0_74542, 
        HIEFFPLA_NET_0_74543, HIEFFPLA_NET_0_74544, 
        HIEFFPLA_NET_0_74545, HIEFFPLA_NET_0_74546, 
        HIEFFPLA_NET_0_74547, HIEFFPLA_NET_0_74548, 
        HIEFFPLA_NET_0_74549, HIEFFPLA_NET_0_74550, 
        HIEFFPLA_NET_0_74551, HIEFFPLA_NET_0_74552, 
        HIEFFPLA_NET_0_74553, HIEFFPLA_NET_0_74554, 
        HIEFFPLA_NET_0_74555, HIEFFPLA_NET_0_74556, 
        HIEFFPLA_NET_0_74557, HIEFFPLA_NET_0_74558, 
        HIEFFPLA_NET_0_74559, HIEFFPLA_NET_0_74560, 
        HIEFFPLA_NET_0_74561, HIEFFPLA_NET_0_74562, 
        HIEFFPLA_NET_0_74563, HIEFFPLA_NET_0_74564, 
        HIEFFPLA_NET_0_74565, HIEFFPLA_NET_0_74566, 
        HIEFFPLA_NET_0_74567, HIEFFPLA_NET_0_74568, 
        HIEFFPLA_NET_0_74569, HIEFFPLA_NET_0_74570, 
        HIEFFPLA_NET_0_74571, HIEFFPLA_NET_0_74572, 
        HIEFFPLA_NET_0_74573, HIEFFPLA_NET_0_74574, 
        HIEFFPLA_NET_0_74575, HIEFFPLA_NET_0_74576, 
        HIEFFPLA_NET_0_74577, HIEFFPLA_NET_0_74578, 
        HIEFFPLA_NET_0_74579, HIEFFPLA_NET_0_74580, 
        HIEFFPLA_NET_0_74581, HIEFFPLA_NET_0_74582, 
        HIEFFPLA_NET_0_74583, HIEFFPLA_NET_0_74584, 
        HIEFFPLA_NET_0_74585, HIEFFPLA_NET_0_74586, 
        HIEFFPLA_NET_0_74587, HIEFFPLA_NET_0_74588, 
        HIEFFPLA_NET_0_74589, HIEFFPLA_NET_0_74590, 
        HIEFFPLA_NET_0_74591, HIEFFPLA_NET_0_74592, 
        HIEFFPLA_NET_0_74593, HIEFFPLA_NET_0_74594, 
        HIEFFPLA_NET_0_74595, HIEFFPLA_NET_0_74596, 
        HIEFFPLA_NET_0_74597, HIEFFPLA_NET_0_74598, 
        HIEFFPLA_NET_0_74599, HIEFFPLA_NET_0_74600, 
        HIEFFPLA_NET_0_74601, HIEFFPLA_NET_0_74602, 
        HIEFFPLA_NET_0_74603, HIEFFPLA_NET_0_74604, 
        HIEFFPLA_NET_0_74605, HIEFFPLA_NET_0_74606, 
        HIEFFPLA_NET_0_74607, HIEFFPLA_NET_0_74608, 
        HIEFFPLA_NET_0_74609, HIEFFPLA_NET_0_74610, 
        HIEFFPLA_NET_0_74611, HIEFFPLA_NET_0_74612, 
        HIEFFPLA_NET_0_74613, HIEFFPLA_NET_0_74614, 
        HIEFFPLA_NET_0_74615, HIEFFPLA_NET_0_74616, 
        HIEFFPLA_NET_0_74617, HIEFFPLA_NET_0_74618, 
        HIEFFPLA_NET_0_74619, HIEFFPLA_NET_0_74620, 
        HIEFFPLA_NET_0_74621, HIEFFPLA_NET_0_74622, 
        HIEFFPLA_NET_0_74623, HIEFFPLA_NET_0_74624, 
        HIEFFPLA_NET_0_74625, HIEFFPLA_NET_0_74626, 
        HIEFFPLA_NET_0_74627, HIEFFPLA_NET_0_74628, 
        HIEFFPLA_NET_0_74629, HIEFFPLA_NET_0_74630, 
        HIEFFPLA_NET_0_74631, HIEFFPLA_NET_0_74632, 
        HIEFFPLA_NET_0_74633, HIEFFPLA_NET_0_74634, 
        HIEFFPLA_NET_0_74635, HIEFFPLA_NET_0_74636, 
        HIEFFPLA_NET_0_74637, HIEFFPLA_NET_0_74638, 
        HIEFFPLA_NET_0_74639, HIEFFPLA_NET_0_74640, 
        HIEFFPLA_NET_0_74641, HIEFFPLA_NET_0_74642, 
        HIEFFPLA_NET_0_74643, HIEFFPLA_NET_0_74644, 
        HIEFFPLA_NET_0_74645, HIEFFPLA_NET_0_74646, 
        HIEFFPLA_NET_0_74647, HIEFFPLA_NET_0_74648, 
        HIEFFPLA_NET_0_74649, HIEFFPLA_NET_0_74650, 
        HIEFFPLA_NET_0_74651, HIEFFPLA_NET_0_74652, 
        HIEFFPLA_NET_0_74653, HIEFFPLA_NET_0_74654, 
        HIEFFPLA_NET_0_74655, HIEFFPLA_NET_0_74656, 
        HIEFFPLA_NET_0_74657, HIEFFPLA_NET_0_74658, 
        HIEFFPLA_NET_0_74659, HIEFFPLA_NET_0_74660, 
        HIEFFPLA_NET_0_74661, HIEFFPLA_NET_0_74662, 
        HIEFFPLA_NET_0_74663, HIEFFPLA_NET_0_74664, 
        HIEFFPLA_NET_0_74665, HIEFFPLA_NET_0_74666, 
        HIEFFPLA_NET_0_74667, HIEFFPLA_NET_0_74668, 
        HIEFFPLA_NET_0_74669, HIEFFPLA_NET_0_74670, 
        HIEFFPLA_NET_0_74671, HIEFFPLA_NET_0_74672, 
        HIEFFPLA_NET_0_74673, HIEFFPLA_NET_0_74674, 
        HIEFFPLA_NET_0_74675, HIEFFPLA_NET_0_74676, 
        HIEFFPLA_NET_0_74677, HIEFFPLA_NET_0_74678, 
        HIEFFPLA_NET_0_74679, HIEFFPLA_NET_0_74680, 
        HIEFFPLA_NET_0_74681, HIEFFPLA_NET_0_74682, 
        HIEFFPLA_NET_0_74683, HIEFFPLA_NET_0_74684, 
        HIEFFPLA_NET_0_74685, HIEFFPLA_NET_0_74686, 
        HIEFFPLA_NET_0_74687, HIEFFPLA_NET_0_74688, 
        HIEFFPLA_NET_0_74689, HIEFFPLA_NET_0_74690, 
        HIEFFPLA_NET_0_74691, HIEFFPLA_NET_0_74692, 
        HIEFFPLA_NET_0_74693, HIEFFPLA_NET_0_74694, 
        HIEFFPLA_NET_0_74695, HIEFFPLA_NET_0_74696, 
        HIEFFPLA_NET_0_74697, HIEFFPLA_NET_0_74698, 
        HIEFFPLA_NET_0_74699, HIEFFPLA_NET_0_74700, 
        HIEFFPLA_NET_0_74701, HIEFFPLA_NET_0_74702, 
        HIEFFPLA_NET_0_74703, HIEFFPLA_NET_0_74704, 
        HIEFFPLA_NET_0_74705, HIEFFPLA_NET_0_74706, 
        HIEFFPLA_NET_0_74707, HIEFFPLA_NET_0_74708, 
        HIEFFPLA_NET_0_74709, HIEFFPLA_NET_0_74710, 
        HIEFFPLA_NET_0_74711, HIEFFPLA_NET_0_74712, 
        HIEFFPLA_NET_0_74713, HIEFFPLA_NET_0_74714, 
        HIEFFPLA_NET_0_74715, HIEFFPLA_NET_0_74716, 
        HIEFFPLA_NET_0_74717, HIEFFPLA_NET_0_74718, 
        HIEFFPLA_NET_0_74719, HIEFFPLA_NET_0_74720, 
        HIEFFPLA_NET_0_74721, HIEFFPLA_NET_0_74722, 
        HIEFFPLA_NET_0_74723, HIEFFPLA_NET_0_74724, 
        HIEFFPLA_NET_0_74725, HIEFFPLA_NET_0_74726, 
        HIEFFPLA_NET_0_74727, HIEFFPLA_NET_0_74728, 
        HIEFFPLA_NET_0_74729, HIEFFPLA_NET_0_74730, 
        HIEFFPLA_NET_0_74731, HIEFFPLA_NET_0_74732, 
        HIEFFPLA_NET_0_74733, HIEFFPLA_NET_0_74734, 
        HIEFFPLA_NET_0_74735, HIEFFPLA_NET_0_74736, 
        HIEFFPLA_NET_0_74737, HIEFFPLA_NET_0_74738, 
        HIEFFPLA_NET_0_74739, HIEFFPLA_NET_0_74740, 
        HIEFFPLA_NET_0_74741, HIEFFPLA_NET_0_74742, 
        HIEFFPLA_NET_0_74743, HIEFFPLA_NET_0_74744, 
        HIEFFPLA_NET_0_74745, HIEFFPLA_NET_0_74746, 
        HIEFFPLA_NET_0_74747, HIEFFPLA_NET_0_74748, 
        HIEFFPLA_NET_0_74749, HIEFFPLA_NET_0_74750, 
        HIEFFPLA_NET_0_74751, HIEFFPLA_NET_0_74752, 
        HIEFFPLA_NET_0_74753, HIEFFPLA_NET_0_74754, 
        HIEFFPLA_NET_0_74755, HIEFFPLA_NET_0_74756, 
        HIEFFPLA_NET_0_74757, HIEFFPLA_NET_0_74758, 
        HIEFFPLA_NET_0_74759, HIEFFPLA_NET_0_74760, 
        HIEFFPLA_NET_0_74761, HIEFFPLA_NET_0_74762, 
        HIEFFPLA_NET_0_74763, HIEFFPLA_NET_0_74764, 
        HIEFFPLA_NET_0_74765, HIEFFPLA_NET_0_74766, 
        HIEFFPLA_NET_0_74767, HIEFFPLA_NET_0_74768, 
        HIEFFPLA_NET_0_74769, HIEFFPLA_NET_0_74770, 
        HIEFFPLA_NET_0_74771, HIEFFPLA_NET_0_74772, 
        HIEFFPLA_NET_0_74773, HIEFFPLA_NET_0_74774, 
        HIEFFPLA_NET_0_74775, HIEFFPLA_NET_0_74776, 
        HIEFFPLA_NET_0_74777, HIEFFPLA_NET_0_74778, 
        HIEFFPLA_NET_0_74779, HIEFFPLA_NET_0_74780, 
        HIEFFPLA_NET_0_74781, HIEFFPLA_NET_0_74782, 
        HIEFFPLA_NET_0_74783, HIEFFPLA_NET_0_74784, 
        HIEFFPLA_NET_0_74785, HIEFFPLA_NET_0_74786, 
        HIEFFPLA_NET_0_74787, HIEFFPLA_NET_0_74788, 
        HIEFFPLA_NET_0_74789, HIEFFPLA_NET_0_74790, 
        HIEFFPLA_NET_0_74791, HIEFFPLA_NET_0_74792, 
        HIEFFPLA_NET_0_74793, HIEFFPLA_NET_0_74794, 
        HIEFFPLA_NET_0_74795, HIEFFPLA_NET_0_74796, 
        HIEFFPLA_NET_0_74797, HIEFFPLA_NET_0_74798, 
        HIEFFPLA_NET_0_74799, HIEFFPLA_NET_0_74800, 
        HIEFFPLA_NET_0_74801, HIEFFPLA_NET_0_74802, 
        HIEFFPLA_NET_0_74803, HIEFFPLA_NET_0_74804, 
        HIEFFPLA_NET_0_74805, HIEFFPLA_NET_0_74806, 
        HIEFFPLA_NET_0_74807, HIEFFPLA_NET_0_74808, 
        HIEFFPLA_NET_0_74809, HIEFFPLA_NET_0_74810, 
        HIEFFPLA_NET_0_74811, HIEFFPLA_NET_0_74812, 
        HIEFFPLA_NET_0_74813, HIEFFPLA_NET_0_74814, 
        HIEFFPLA_NET_0_74815, HIEFFPLA_NET_0_74816, 
        HIEFFPLA_NET_0_74817, HIEFFPLA_NET_0_74818, 
        HIEFFPLA_NET_0_74819, HIEFFPLA_NET_0_74820, 
        HIEFFPLA_NET_0_74821, HIEFFPLA_NET_0_74822, 
        HIEFFPLA_NET_0_74823, HIEFFPLA_NET_0_74824, 
        HIEFFPLA_NET_0_74825, HIEFFPLA_NET_0_74826, 
        HIEFFPLA_NET_0_74827, HIEFFPLA_NET_0_74828, 
        HIEFFPLA_NET_0_74829, HIEFFPLA_NET_0_74830, 
        HIEFFPLA_NET_0_74831, HIEFFPLA_NET_0_74832, 
        HIEFFPLA_NET_0_74833, HIEFFPLA_NET_0_74834, 
        HIEFFPLA_NET_0_74835, HIEFFPLA_NET_0_74836, 
        HIEFFPLA_NET_0_74837, HIEFFPLA_NET_0_74838, 
        HIEFFPLA_NET_0_74839, HIEFFPLA_NET_0_74840, 
        HIEFFPLA_NET_0_74841, HIEFFPLA_NET_0_74842, 
        HIEFFPLA_NET_0_74843, HIEFFPLA_NET_0_74844, 
        HIEFFPLA_NET_0_74845, HIEFFPLA_NET_0_74846, 
        HIEFFPLA_NET_0_74847, HIEFFPLA_NET_0_74848, 
        HIEFFPLA_NET_0_74849, HIEFFPLA_NET_0_74850, 
        HIEFFPLA_NET_0_74851, HIEFFPLA_NET_0_74852, 
        HIEFFPLA_NET_0_74853, HIEFFPLA_NET_0_74854, 
        HIEFFPLA_NET_0_74855, HIEFFPLA_NET_0_74856, 
        HIEFFPLA_NET_0_74857, HIEFFPLA_NET_0_74858, 
        HIEFFPLA_NET_0_74859, HIEFFPLA_NET_0_74860, 
        HIEFFPLA_NET_0_74861, HIEFFPLA_NET_0_74862, 
        HIEFFPLA_NET_0_74863, HIEFFPLA_NET_0_74864, 
        HIEFFPLA_NET_0_74865, HIEFFPLA_NET_0_74866, 
        HIEFFPLA_NET_0_74867, HIEFFPLA_NET_0_74868, 
        HIEFFPLA_NET_0_74869, HIEFFPLA_NET_0_74870, 
        HIEFFPLA_NET_0_74871, HIEFFPLA_NET_0_74872, 
        HIEFFPLA_NET_0_74873, HIEFFPLA_NET_0_74874, 
        HIEFFPLA_NET_0_74875, HIEFFPLA_NET_0_74876, 
        HIEFFPLA_NET_0_74877, HIEFFPLA_NET_0_74878, 
        HIEFFPLA_NET_0_74879, HIEFFPLA_NET_0_74880, 
        HIEFFPLA_NET_0_74881, HIEFFPLA_NET_0_74882, 
        HIEFFPLA_NET_0_74883, HIEFFPLA_NET_0_74884, 
        HIEFFPLA_NET_0_74885, HIEFFPLA_NET_0_74886, 
        HIEFFPLA_NET_0_74887, HIEFFPLA_NET_0_74888, 
        HIEFFPLA_NET_0_74889, HIEFFPLA_NET_0_74890, 
        HIEFFPLA_NET_0_74891, HIEFFPLA_NET_0_74892, 
        HIEFFPLA_NET_0_74893, HIEFFPLA_NET_0_74894, 
        HIEFFPLA_NET_0_74895, HIEFFPLA_NET_0_74896, 
        HIEFFPLA_NET_0_74897, HIEFFPLA_NET_0_74898, 
        HIEFFPLA_NET_0_74899, HIEFFPLA_NET_0_74900, 
        HIEFFPLA_NET_0_74901, HIEFFPLA_NET_0_74902, 
        HIEFFPLA_NET_0_74903, HIEFFPLA_NET_0_74904, 
        HIEFFPLA_NET_0_74905, HIEFFPLA_NET_0_74906, 
        HIEFFPLA_NET_0_74907, HIEFFPLA_NET_0_74908, 
        HIEFFPLA_NET_0_74909, HIEFFPLA_NET_0_74910, 
        HIEFFPLA_NET_0_74911, HIEFFPLA_NET_0_74912, 
        HIEFFPLA_NET_0_74913, HIEFFPLA_NET_0_74914, 
        HIEFFPLA_NET_0_74915, HIEFFPLA_NET_0_74916, 
        HIEFFPLA_NET_0_74917, HIEFFPLA_NET_0_74918, 
        HIEFFPLA_NET_0_74919, HIEFFPLA_NET_0_74920, 
        HIEFFPLA_NET_0_74921, HIEFFPLA_NET_0_74922, 
        HIEFFPLA_NET_0_74923, HIEFFPLA_NET_0_74924, 
        HIEFFPLA_NET_0_74925, HIEFFPLA_NET_0_74926, 
        HIEFFPLA_NET_0_74927, HIEFFPLA_NET_0_74928, 
        HIEFFPLA_NET_0_74929, HIEFFPLA_NET_0_74930, 
        HIEFFPLA_NET_0_74931, HIEFFPLA_NET_0_74932, 
        HIEFFPLA_NET_0_74933, HIEFFPLA_NET_0_74934, 
        HIEFFPLA_NET_0_74935, HIEFFPLA_NET_0_74936, 
        HIEFFPLA_NET_0_74937, HIEFFPLA_NET_0_74938, 
        HIEFFPLA_NET_0_74939, HIEFFPLA_NET_0_74940, 
        HIEFFPLA_NET_0_74941, HIEFFPLA_NET_0_74942, 
        HIEFFPLA_NET_0_74943, HIEFFPLA_NET_0_74944, 
        HIEFFPLA_NET_0_74945, HIEFFPLA_NET_0_74946, 
        HIEFFPLA_NET_0_74947, HIEFFPLA_NET_0_74948, 
        HIEFFPLA_NET_0_74949, HIEFFPLA_NET_0_74950, 
        HIEFFPLA_NET_0_74951, HIEFFPLA_NET_0_74952, 
        HIEFFPLA_NET_0_74953, HIEFFPLA_NET_0_74954, 
        HIEFFPLA_NET_0_74955, HIEFFPLA_NET_0_74956, 
        HIEFFPLA_NET_0_74957, HIEFFPLA_NET_0_74958, 
        HIEFFPLA_NET_0_74959, HIEFFPLA_NET_0_74960, 
        HIEFFPLA_NET_0_74961, HIEFFPLA_NET_0_74962, 
        HIEFFPLA_NET_0_74963, HIEFFPLA_NET_0_74964, 
        HIEFFPLA_NET_0_74965, HIEFFPLA_NET_0_74966, 
        HIEFFPLA_NET_0_74967, HIEFFPLA_NET_0_74968, 
        HIEFFPLA_NET_0_74969, HIEFFPLA_NET_0_74970, 
        HIEFFPLA_NET_0_74971, HIEFFPLA_NET_0_74972, 
        HIEFFPLA_NET_0_74973, HIEFFPLA_NET_0_74974, 
        HIEFFPLA_NET_0_74975, HIEFFPLA_NET_0_74976, 
        HIEFFPLA_NET_0_74977, HIEFFPLA_NET_0_74978, 
        HIEFFPLA_NET_0_74979, HIEFFPLA_NET_0_74980, 
        HIEFFPLA_NET_0_74981, HIEFFPLA_NET_0_74982, 
        HIEFFPLA_NET_0_74983, HIEFFPLA_NET_0_74984, 
        HIEFFPLA_NET_0_74985, HIEFFPLA_NET_0_74986, 
        HIEFFPLA_NET_0_74987, HIEFFPLA_NET_0_74988, 
        HIEFFPLA_NET_0_74989, HIEFFPLA_NET_0_74990, 
        HIEFFPLA_NET_0_74991, HIEFFPLA_NET_0_74992, 
        HIEFFPLA_NET_0_74993, HIEFFPLA_NET_0_74994, 
        HIEFFPLA_NET_0_74995, HIEFFPLA_NET_0_74996, 
        HIEFFPLA_NET_0_74997, HIEFFPLA_NET_0_74998, 
        HIEFFPLA_NET_0_74999, HIEFFPLA_NET_0_75000, 
        HIEFFPLA_NET_0_75001, HIEFFPLA_NET_0_75002, 
        HIEFFPLA_NET_0_75003, HIEFFPLA_NET_0_75004, 
        HIEFFPLA_NET_0_75005, HIEFFPLA_NET_0_75006, 
        HIEFFPLA_NET_0_75007, HIEFFPLA_NET_0_75008, 
        HIEFFPLA_NET_0_75009, HIEFFPLA_NET_0_75010, 
        HIEFFPLA_NET_0_75011, HIEFFPLA_NET_0_75012, 
        HIEFFPLA_NET_0_75013, HIEFFPLA_NET_0_75014, 
        HIEFFPLA_NET_0_75015, HIEFFPLA_NET_0_75016, 
        HIEFFPLA_NET_0_75017, HIEFFPLA_NET_0_75018, 
        HIEFFPLA_NET_0_75019, HIEFFPLA_NET_0_75020, 
        HIEFFPLA_NET_0_75021, HIEFFPLA_NET_0_75022, 
        HIEFFPLA_NET_0_75023, HIEFFPLA_NET_0_75024, 
        HIEFFPLA_NET_0_75025, HIEFFPLA_NET_0_75026, 
        HIEFFPLA_NET_0_75027, HIEFFPLA_NET_0_75028, 
        HIEFFPLA_NET_0_75029, HIEFFPLA_NET_0_75030, 
        HIEFFPLA_NET_0_75031, HIEFFPLA_NET_0_75032, 
        HIEFFPLA_NET_0_75033, HIEFFPLA_NET_0_75034, 
        HIEFFPLA_NET_0_75035, HIEFFPLA_NET_0_75036, 
        HIEFFPLA_NET_0_75037, HIEFFPLA_NET_0_75038, 
        HIEFFPLA_NET_0_75039, HIEFFPLA_NET_0_75040, 
        HIEFFPLA_NET_0_75041, HIEFFPLA_NET_0_75042, 
        HIEFFPLA_NET_0_75043, HIEFFPLA_NET_0_75044, 
        HIEFFPLA_NET_0_75045, HIEFFPLA_NET_0_75046, 
        HIEFFPLA_NET_0_75047, HIEFFPLA_NET_0_75048, 
        HIEFFPLA_NET_0_75049, HIEFFPLA_NET_0_75050, 
        HIEFFPLA_NET_0_75051, HIEFFPLA_NET_0_75052, 
        HIEFFPLA_NET_0_75053, HIEFFPLA_NET_0_75054, 
        HIEFFPLA_NET_0_75055, HIEFFPLA_NET_0_75056, 
        HIEFFPLA_NET_0_75057, HIEFFPLA_NET_0_75058, 
        HIEFFPLA_NET_0_75059, HIEFFPLA_NET_0_75060, 
        HIEFFPLA_NET_0_75061, HIEFFPLA_NET_0_75062, 
        HIEFFPLA_NET_0_75063, HIEFFPLA_NET_0_75064, 
        HIEFFPLA_NET_0_75065, HIEFFPLA_NET_0_75066, 
        HIEFFPLA_NET_0_75067, HIEFFPLA_NET_0_75068, 
        HIEFFPLA_NET_0_75069, HIEFFPLA_NET_0_75070, 
        HIEFFPLA_NET_0_75071, HIEFFPLA_NET_0_75072, 
        HIEFFPLA_NET_0_75073, HIEFFPLA_NET_0_75074, 
        HIEFFPLA_NET_0_75075, HIEFFPLA_NET_0_75076, 
        HIEFFPLA_NET_0_75077, HIEFFPLA_NET_0_75078, 
        HIEFFPLA_NET_0_75079, HIEFFPLA_NET_0_75080, 
        HIEFFPLA_NET_0_75081, HIEFFPLA_NET_0_75082, 
        HIEFFPLA_NET_0_75083, HIEFFPLA_NET_0_75084, 
        HIEFFPLA_NET_0_75085, HIEFFPLA_NET_0_75086, 
        HIEFFPLA_NET_0_75087, HIEFFPLA_NET_0_75088, 
        HIEFFPLA_NET_0_75089, HIEFFPLA_NET_0_75090, 
        HIEFFPLA_NET_0_75091, HIEFFPLA_NET_0_75092, 
        HIEFFPLA_NET_0_75093, HIEFFPLA_NET_0_75094, 
        HIEFFPLA_NET_0_75095, HIEFFPLA_NET_0_75096, 
        HIEFFPLA_NET_0_75097, HIEFFPLA_NET_0_75098, 
        HIEFFPLA_NET_0_75099, HIEFFPLA_NET_0_75100, 
        HIEFFPLA_NET_0_75101, HIEFFPLA_NET_0_75102, 
        HIEFFPLA_NET_0_75103, HIEFFPLA_NET_0_75104, 
        HIEFFPLA_NET_0_75105, HIEFFPLA_NET_0_75106, 
        HIEFFPLA_NET_0_75107, HIEFFPLA_NET_0_75108, 
        HIEFFPLA_NET_0_75109, HIEFFPLA_NET_0_75110, 
        HIEFFPLA_NET_0_75111, HIEFFPLA_NET_0_75112, 
        HIEFFPLA_NET_0_75113, HIEFFPLA_NET_0_75114, 
        HIEFFPLA_NET_0_75115, HIEFFPLA_NET_0_75116, 
        HIEFFPLA_NET_0_75117, HIEFFPLA_NET_0_75118, 
        HIEFFPLA_NET_0_75119, HIEFFPLA_NET_0_75120, 
        HIEFFPLA_NET_0_75121, HIEFFPLA_NET_0_75122, 
        HIEFFPLA_NET_0_75123, HIEFFPLA_NET_0_75124, 
        HIEFFPLA_NET_0_75125, HIEFFPLA_NET_0_75126, 
        HIEFFPLA_NET_0_75127, HIEFFPLA_NET_0_75128, 
        HIEFFPLA_NET_0_75129, HIEFFPLA_NET_0_75130, 
        HIEFFPLA_NET_0_75131, HIEFFPLA_NET_0_75132, 
        HIEFFPLA_NET_0_75133, HIEFFPLA_NET_0_75134, 
        HIEFFPLA_NET_0_75135, HIEFFPLA_NET_0_75136, 
        HIEFFPLA_NET_0_75137, HIEFFPLA_NET_0_75138, 
        HIEFFPLA_NET_0_75139, HIEFFPLA_NET_0_75140, 
        HIEFFPLA_NET_0_75141, HIEFFPLA_NET_0_75142, 
        HIEFFPLA_NET_0_75143, HIEFFPLA_NET_0_75144, 
        HIEFFPLA_NET_0_75145, HIEFFPLA_NET_0_75146, 
        HIEFFPLA_NET_0_75147, HIEFFPLA_NET_0_75148, 
        HIEFFPLA_NET_0_75149, HIEFFPLA_NET_0_75150, 
        HIEFFPLA_NET_0_75151, HIEFFPLA_NET_0_75152, 
        HIEFFPLA_NET_0_75153, HIEFFPLA_NET_0_75154, 
        HIEFFPLA_NET_0_75155, HIEFFPLA_NET_0_75156, 
        HIEFFPLA_NET_0_75157, HIEFFPLA_NET_0_75158, 
        HIEFFPLA_NET_0_75159, HIEFFPLA_NET_0_75160, 
        HIEFFPLA_NET_0_75161, HIEFFPLA_NET_0_75162, 
        HIEFFPLA_NET_0_75163, HIEFFPLA_NET_0_75164, 
        HIEFFPLA_NET_0_75165, HIEFFPLA_NET_0_75166, 
        HIEFFPLA_NET_0_75167, HIEFFPLA_NET_0_75168, 
        HIEFFPLA_NET_0_75169, HIEFFPLA_NET_0_75170, 
        HIEFFPLA_NET_0_75171, HIEFFPLA_NET_0_75172, 
        HIEFFPLA_NET_0_75173, HIEFFPLA_NET_0_75174, 
        HIEFFPLA_NET_0_75175, HIEFFPLA_NET_0_75176, 
        HIEFFPLA_NET_0_75177, HIEFFPLA_NET_0_75178, 
        HIEFFPLA_NET_0_75179, HIEFFPLA_NET_0_75180, 
        HIEFFPLA_NET_0_75181, HIEFFPLA_NET_0_75182, 
        HIEFFPLA_NET_0_75183, HIEFFPLA_NET_0_75184, 
        HIEFFPLA_NET_0_75185, HIEFFPLA_NET_0_75186, 
        HIEFFPLA_NET_0_75187, HIEFFPLA_NET_0_75188, 
        HIEFFPLA_NET_0_75189, HIEFFPLA_NET_0_75190, 
        HIEFFPLA_NET_0_75191, HIEFFPLA_NET_0_75192, 
        HIEFFPLA_NET_0_75193, HIEFFPLA_NET_0_75194, 
        HIEFFPLA_NET_0_75195, HIEFFPLA_NET_0_75196, 
        HIEFFPLA_NET_0_75197, HIEFFPLA_NET_0_75198, 
        HIEFFPLA_NET_0_75199, HIEFFPLA_NET_0_75200, 
        HIEFFPLA_NET_0_75201, HIEFFPLA_NET_0_75202, 
        HIEFFPLA_NET_0_75203, HIEFFPLA_NET_0_75204, 
        HIEFFPLA_NET_0_75205, HIEFFPLA_NET_0_75206, 
        HIEFFPLA_NET_0_75207, HIEFFPLA_NET_0_75208, 
        HIEFFPLA_NET_0_75209, HIEFFPLA_NET_0_75210, 
        HIEFFPLA_NET_0_75211, HIEFFPLA_NET_0_75212, 
        HIEFFPLA_NET_0_75213, HIEFFPLA_NET_0_75214, 
        HIEFFPLA_NET_0_75215, HIEFFPLA_NET_0_75216, 
        HIEFFPLA_NET_0_75217, HIEFFPLA_NET_0_75218, 
        HIEFFPLA_NET_0_75219, HIEFFPLA_NET_0_75220, 
        HIEFFPLA_NET_0_75221, HIEFFPLA_NET_0_75222, 
        HIEFFPLA_NET_0_75223, HIEFFPLA_NET_0_75224, 
        HIEFFPLA_NET_0_75225, HIEFFPLA_NET_0_75226, 
        HIEFFPLA_NET_0_75227, HIEFFPLA_NET_0_75228, 
        HIEFFPLA_NET_0_75229, HIEFFPLA_NET_0_75230, 
        HIEFFPLA_NET_0_75231, HIEFFPLA_NET_0_75232, 
        HIEFFPLA_NET_0_75233, HIEFFPLA_NET_0_75234, 
        HIEFFPLA_NET_0_75235, HIEFFPLA_NET_0_75236, 
        HIEFFPLA_NET_0_75237, HIEFFPLA_NET_0_75238, 
        HIEFFPLA_NET_0_75239, HIEFFPLA_NET_0_75240, 
        HIEFFPLA_NET_0_75241, HIEFFPLA_NET_0_75242, 
        HIEFFPLA_NET_0_75243, HIEFFPLA_NET_0_75244, 
        HIEFFPLA_NET_0_75245, HIEFFPLA_NET_0_75246, 
        HIEFFPLA_NET_0_75247, HIEFFPLA_NET_0_75248, 
        HIEFFPLA_NET_0_75249, HIEFFPLA_NET_0_75250, 
        HIEFFPLA_NET_0_75251, HIEFFPLA_NET_0_75252, 
        HIEFFPLA_NET_0_75253, HIEFFPLA_NET_0_75254, 
        HIEFFPLA_NET_0_75255, HIEFFPLA_NET_0_75256, 
        HIEFFPLA_NET_0_75257, HIEFFPLA_NET_0_75258, 
        HIEFFPLA_NET_0_75259, HIEFFPLA_NET_0_75260, 
        HIEFFPLA_NET_0_75261, HIEFFPLA_NET_0_75262, 
        HIEFFPLA_NET_0_75263, HIEFFPLA_NET_0_75264, 
        HIEFFPLA_NET_0_75265, HIEFFPLA_NET_0_75266, 
        HIEFFPLA_NET_0_75267, HIEFFPLA_NET_0_75268, 
        HIEFFPLA_NET_0_75269, HIEFFPLA_NET_0_75270, 
        HIEFFPLA_NET_0_75271, HIEFFPLA_NET_0_75272, 
        HIEFFPLA_NET_0_75273, HIEFFPLA_NET_0_75274, 
        HIEFFPLA_NET_0_75275, HIEFFPLA_NET_0_75276, 
        HIEFFPLA_NET_0_75277, HIEFFPLA_NET_0_75278, 
        HIEFFPLA_NET_0_75279, HIEFFPLA_NET_0_75280, 
        HIEFFPLA_NET_0_75281, HIEFFPLA_NET_0_75282, 
        HIEFFPLA_NET_0_75283, HIEFFPLA_NET_0_75284, 
        HIEFFPLA_NET_0_75285, HIEFFPLA_NET_0_75286, 
        HIEFFPLA_NET_0_75287, HIEFFPLA_NET_0_75288, 
        HIEFFPLA_NET_0_75289, HIEFFPLA_NET_0_75290, 
        HIEFFPLA_NET_0_75291, HIEFFPLA_NET_0_75292, 
        HIEFFPLA_NET_0_75293, HIEFFPLA_NET_0_75294, 
        HIEFFPLA_NET_0_75295, HIEFFPLA_NET_0_75296, 
        HIEFFPLA_NET_0_75297, HIEFFPLA_NET_0_75298, 
        HIEFFPLA_NET_0_75299, HIEFFPLA_NET_0_75300, 
        HIEFFPLA_NET_0_75301, HIEFFPLA_NET_0_75302, 
        HIEFFPLA_NET_0_75303, HIEFFPLA_NET_0_75304, 
        HIEFFPLA_NET_0_75305, HIEFFPLA_NET_0_75306, 
        HIEFFPLA_NET_0_75307, HIEFFPLA_NET_0_75308, 
        HIEFFPLA_NET_0_75309, HIEFFPLA_NET_0_75310, 
        HIEFFPLA_NET_0_75311, HIEFFPLA_NET_0_75312, 
        HIEFFPLA_NET_0_75313, HIEFFPLA_NET_0_75314, 
        HIEFFPLA_NET_0_75315, HIEFFPLA_NET_0_75316, 
        HIEFFPLA_NET_0_75317, HIEFFPLA_NET_0_75318, 
        HIEFFPLA_NET_0_75319, HIEFFPLA_NET_0_75320, 
        HIEFFPLA_NET_0_75321, HIEFFPLA_NET_0_75322, 
        HIEFFPLA_NET_0_75323, HIEFFPLA_NET_0_75324, 
        HIEFFPLA_NET_0_75325, HIEFFPLA_NET_0_75326, 
        HIEFFPLA_NET_0_75327, HIEFFPLA_NET_0_75328, 
        HIEFFPLA_NET_0_75329, HIEFFPLA_NET_0_75330, 
        HIEFFPLA_NET_0_75331, HIEFFPLA_NET_0_75336, 
        HIEFFPLA_NET_0_75338, HIEFFPLA_NET_0_75339, 
        HIEFFPLA_NET_0_75340, HIEFFPLA_NET_0_75341, 
        HIEFFPLA_NET_0_75343, HIEFFPLA_NET_0_75344, 
        HIEFFPLA_NET_0_75345, HIEFFPLA_NET_0_75346, 
        HIEFFPLA_NET_0_75347, HIEFFPLA_NET_0_75348, 
        HIEFFPLA_NET_0_75349, HIEFFPLA_NET_0_75350, 
        HIEFFPLA_NET_0_75351, HIEFFPLA_NET_0_75352, 
        HIEFFPLA_NET_0_75353, HIEFFPLA_NET_0_75354, 
        HIEFFPLA_NET_0_75355, HIEFFPLA_NET_0_75356, 
        HIEFFPLA_NET_0_75357, HIEFFPLA_NET_0_75358, 
        HIEFFPLA_NET_0_75359, HIEFFPLA_NET_0_75360, 
        HIEFFPLA_NET_0_75361, HIEFFPLA_NET_0_75362, 
        HIEFFPLA_NET_0_75363, HIEFFPLA_NET_0_75364, 
        HIEFFPLA_NET_0_75366, HIEFFPLA_NET_0_75367, 
        HIEFFPLA_NET_0_75368, HIEFFPLA_NET_0_75369, 
        HIEFFPLA_NET_0_75370, HIEFFPLA_NET_0_75371, 
        HIEFFPLA_NET_0_75372, HIEFFPLA_NET_0_75373, 
        HIEFFPLA_NET_0_75374, HIEFFPLA_NET_0_75375, 
        HIEFFPLA_NET_0_75376, HIEFFPLA_NET_0_75378, 
        HIEFFPLA_NET_0_75380, HIEFFPLA_NET_0_75381, 
        HIEFFPLA_NET_0_75382, HIEFFPLA_NET_0_75383, 
        HIEFFPLA_NET_0_75384, HIEFFPLA_NET_0_75385, 
        HIEFFPLA_NET_0_75386, HIEFFPLA_NET_0_75387, 
        HIEFFPLA_NET_0_75388, HIEFFPLA_NET_0_75389, 
        HIEFFPLA_NET_0_75390, HIEFFPLA_NET_0_75391, 
        HIEFFPLA_NET_0_75392, HIEFFPLA_NET_0_75393, 
        HIEFFPLA_NET_0_75394, HIEFFPLA_NET_0_75395, 
        HIEFFPLA_NET_0_75396, HIEFFPLA_NET_0_75397, 
        HIEFFPLA_NET_0_75398, HIEFFPLA_NET_0_75399, 
        HIEFFPLA_NET_0_75400, HIEFFPLA_NET_0_75401, 
        HIEFFPLA_NET_0_75402, HIEFFPLA_NET_0_75403, 
        HIEFFPLA_NET_0_75404, HIEFFPLA_NET_0_75405, 
        HIEFFPLA_NET_0_75406, HIEFFPLA_NET_0_75407, 
        HIEFFPLA_NET_0_75408, HIEFFPLA_NET_0_75409, 
        HIEFFPLA_NET_0_75410, HIEFFPLA_NET_0_75411, 
        HIEFFPLA_NET_0_75412, HIEFFPLA_NET_0_75413, 
        HIEFFPLA_NET_0_75414, HIEFFPLA_NET_0_75415, 
        HIEFFPLA_NET_0_75416, HIEFFPLA_NET_0_75417, 
        HIEFFPLA_NET_0_75418, HIEFFPLA_NET_0_75419, 
        HIEFFPLA_NET_0_75420, HIEFFPLA_NET_0_75421, 
        HIEFFPLA_NET_0_75422, HIEFFPLA_NET_0_75423, 
        HIEFFPLA_NET_0_75424, HIEFFPLA_NET_0_75425, 
        HIEFFPLA_NET_0_75426, HIEFFPLA_NET_0_75427, 
        HIEFFPLA_NET_0_75428, HIEFFPLA_NET_0_75429, 
        HIEFFPLA_NET_0_75430, HIEFFPLA_NET_0_75431, 
        HIEFFPLA_NET_0_75432, HIEFFPLA_NET_0_75433, 
        HIEFFPLA_NET_0_75434, HIEFFPLA_NET_0_75435, 
        HIEFFPLA_NET_0_75436, HIEFFPLA_NET_0_75437, 
        HIEFFPLA_NET_0_75438, HIEFFPLA_NET_0_75439, 
        HIEFFPLA_NET_0_75440, HIEFFPLA_NET_0_75441, 
        HIEFFPLA_NET_0_75442, HIEFFPLA_NET_0_75443, 
        HIEFFPLA_NET_0_75444, HIEFFPLA_NET_0_75445, 
        HIEFFPLA_NET_0_75446, HIEFFPLA_NET_0_75447, 
        HIEFFPLA_NET_0_75448, HIEFFPLA_NET_0_75449, 
        HIEFFPLA_NET_0_75450, HIEFFPLA_NET_0_75451, 
        HIEFFPLA_NET_0_75452, HIEFFPLA_NET_0_75453, 
        HIEFFPLA_NET_0_75454, HIEFFPLA_NET_0_75455, 
        HIEFFPLA_NET_0_75456, HIEFFPLA_NET_0_75457, 
        HIEFFPLA_NET_0_75458, HIEFFPLA_NET_0_75459, 
        HIEFFPLA_NET_0_75460, HIEFFPLA_NET_0_75461, 
        HIEFFPLA_NET_0_75462, HIEFFPLA_NET_0_75463, 
        HIEFFPLA_NET_0_75464, HIEFFPLA_NET_0_75465, 
        HIEFFPLA_NET_0_75466, HIEFFPLA_NET_0_75467, 
        HIEFFPLA_NET_0_75468, HIEFFPLA_NET_0_75469, 
        HIEFFPLA_NET_0_75470, HIEFFPLA_NET_0_75471, 
        HIEFFPLA_NET_0_75472, HIEFFPLA_NET_0_75473, 
        HIEFFPLA_NET_0_75474, HIEFFPLA_NET_0_75475, 
        HIEFFPLA_NET_0_75476, HIEFFPLA_NET_0_75477, 
        HIEFFPLA_NET_0_75478, HIEFFPLA_NET_0_75479, 
        HIEFFPLA_NET_0_75480, HIEFFPLA_NET_0_75481, 
        HIEFFPLA_NET_0_75482, HIEFFPLA_NET_0_75483, 
        HIEFFPLA_NET_0_75484, HIEFFPLA_NET_0_75485, 
        HIEFFPLA_NET_0_75486, HIEFFPLA_NET_0_75487, 
        HIEFFPLA_NET_0_75488, HIEFFPLA_NET_0_75489, 
        HIEFFPLA_NET_0_75490, HIEFFPLA_NET_0_75491, 
        HIEFFPLA_NET_0_75492, HIEFFPLA_NET_0_75493, 
        HIEFFPLA_NET_0_75494, HIEFFPLA_NET_0_75495, 
        HIEFFPLA_NET_0_75496, HIEFFPLA_NET_0_75497, 
        HIEFFPLA_NET_0_75498, HIEFFPLA_NET_0_75499, 
        HIEFFPLA_NET_0_75500, HIEFFPLA_NET_0_75501, 
        HIEFFPLA_NET_0_75502, HIEFFPLA_NET_0_75503, 
        HIEFFPLA_NET_0_75504, HIEFFPLA_NET_0_75505, 
        HIEFFPLA_NET_0_75506, HIEFFPLA_NET_0_75507, 
        HIEFFPLA_NET_0_75508, HIEFFPLA_NET_0_75509, 
        HIEFFPLA_NET_0_75510, HIEFFPLA_NET_0_75511, 
        HIEFFPLA_NET_0_75512, HIEFFPLA_NET_0_75513, 
        HIEFFPLA_NET_0_75514, HIEFFPLA_NET_0_75515, 
        HIEFFPLA_NET_0_75516, HIEFFPLA_NET_0_75517, 
        HIEFFPLA_NET_0_75518, HIEFFPLA_NET_0_75519, 
        HIEFFPLA_NET_0_75520, HIEFFPLA_NET_0_75521, 
        HIEFFPLA_NET_0_75522, HIEFFPLA_NET_0_75523, 
        HIEFFPLA_NET_0_75524, HIEFFPLA_NET_0_75525, 
        HIEFFPLA_NET_0_75526, HIEFFPLA_NET_0_75527, 
        HIEFFPLA_NET_0_75528, HIEFFPLA_NET_0_75529, 
        HIEFFPLA_NET_0_75530, HIEFFPLA_NET_0_75531, 
        HIEFFPLA_NET_0_75532, HIEFFPLA_NET_0_75533, 
        HIEFFPLA_NET_0_75534, HIEFFPLA_NET_0_75535, 
        HIEFFPLA_NET_0_75536, HIEFFPLA_NET_0_75537, 
        HIEFFPLA_NET_0_75538, HIEFFPLA_NET_0_75539, 
        HIEFFPLA_NET_0_75540, HIEFFPLA_NET_0_75541, 
        HIEFFPLA_NET_0_75542, HIEFFPLA_NET_0_75543, 
        HIEFFPLA_NET_0_75544, HIEFFPLA_NET_0_75545, 
        HIEFFPLA_NET_0_75546, HIEFFPLA_NET_0_75547, 
        HIEFFPLA_NET_0_75548, HIEFFPLA_NET_0_75549, 
        HIEFFPLA_NET_0_75550, HIEFFPLA_NET_0_75551, 
        HIEFFPLA_NET_0_75552, HIEFFPLA_NET_0_75553, 
        HIEFFPLA_NET_0_75554, HIEFFPLA_NET_0_75555, 
        HIEFFPLA_NET_0_75556, HIEFFPLA_NET_0_75557, 
        HIEFFPLA_NET_0_75558, HIEFFPLA_NET_0_75559, 
        HIEFFPLA_NET_0_75560, HIEFFPLA_NET_0_75561, 
        HIEFFPLA_NET_0_75562, HIEFFPLA_NET_0_75563, 
        HIEFFPLA_NET_0_75564, HIEFFPLA_NET_0_75565, 
        HIEFFPLA_NET_0_75566, HIEFFPLA_NET_0_75567, 
        HIEFFPLA_NET_0_75568, HIEFFPLA_NET_0_75569, 
        HIEFFPLA_NET_0_75570, HIEFFPLA_NET_0_75571, 
        HIEFFPLA_NET_0_75572, HIEFFPLA_NET_0_75573, 
        HIEFFPLA_NET_0_75574, HIEFFPLA_NET_0_75575, 
        HIEFFPLA_NET_0_75576, HIEFFPLA_NET_0_75577, 
        HIEFFPLA_NET_0_75578, HIEFFPLA_NET_0_75579, 
        HIEFFPLA_NET_0_75580, HIEFFPLA_NET_0_75581, 
        HIEFFPLA_NET_0_75582, HIEFFPLA_NET_0_75583, 
        HIEFFPLA_NET_0_75584, HIEFFPLA_NET_0_75585, 
        HIEFFPLA_NET_0_75586, HIEFFPLA_NET_0_75587, 
        HIEFFPLA_NET_0_75588, HIEFFPLA_NET_0_75589, 
        HIEFFPLA_NET_0_75590, HIEFFPLA_NET_0_75591, 
        HIEFFPLA_NET_0_75592, HIEFFPLA_NET_0_75593, 
        HIEFFPLA_NET_0_75594, HIEFFPLA_NET_0_75595, 
        HIEFFPLA_NET_0_75596, HIEFFPLA_NET_0_75597, 
        HIEFFPLA_NET_0_75598, HIEFFPLA_NET_0_75599, 
        HIEFFPLA_NET_0_75600, HIEFFPLA_NET_0_75601, 
        HIEFFPLA_NET_0_75602, HIEFFPLA_NET_0_75603, 
        HIEFFPLA_NET_0_75604, HIEFFPLA_NET_0_75605, 
        HIEFFPLA_NET_0_75606, HIEFFPLA_NET_0_75607, 
        HIEFFPLA_NET_0_75608, HIEFFPLA_NET_0_75609, 
        HIEFFPLA_NET_0_75610, HIEFFPLA_NET_0_75611, 
        HIEFFPLA_NET_0_75612, HIEFFPLA_NET_0_75613, 
        HIEFFPLA_NET_0_75614, HIEFFPLA_NET_0_75615, 
        HIEFFPLA_NET_0_75616, HIEFFPLA_NET_0_75617, 
        HIEFFPLA_NET_0_75618, HIEFFPLA_NET_0_75619, 
        HIEFFPLA_NET_0_75620, HIEFFPLA_NET_0_75621, 
        HIEFFPLA_NET_0_75622, HIEFFPLA_NET_0_75623, 
        HIEFFPLA_NET_0_75624, HIEFFPLA_NET_0_75625, 
        HIEFFPLA_NET_0_75626, HIEFFPLA_NET_0_75627, 
        HIEFFPLA_NET_0_75628, HIEFFPLA_NET_0_75629, 
        HIEFFPLA_NET_0_75630, HIEFFPLA_NET_0_75631, 
        HIEFFPLA_NET_0_75632, HIEFFPLA_NET_0_75633, 
        HIEFFPLA_NET_0_75634, HIEFFPLA_NET_0_75635, 
        HIEFFPLA_NET_0_75636, HIEFFPLA_NET_0_75637, 
        HIEFFPLA_NET_0_75638, HIEFFPLA_NET_0_88380, 
        HIEFFPLA_NET_0_88381, HIEFFPLA_NET_0_88382, 
        HIEFFPLA_NET_0_88383, HIEFFPLA_NET_0_88384, 
        HIEFFPLA_NET_0_88385, HIEFFPLA_NET_0_88386, 
        HIEFFPLA_NET_0_88387, HIEFFPLA_NET_0_89694, 
        HIEFFPLA_NET_0_89700, HIEFFPLA_NET_0_89701, 
        \I2C_PassThrough_0/cnt[0]_net_1\, 
        \I2C_PassThrough_0/cnt[1]_net_1\, 
        \I2C_PassThrough_0/cnt[2]_net_1\, 
        \I2C_PassThrough_0/cnt[3]_net_1\, 
        \I2C_PassThrough_0/cnt[4]_net_1\, 
        \I2C_PassThrough_0/state[0]_net_1\, 
        \I2C_PassThrough_0/state[1]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[0]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[1]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[2]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[3]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[4]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[5]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[6]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[7]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[8]_net_1\, 
        \Pressure_Signal_Debounce_0/ms_cnt[9]_net_1\, 
        \Pressure_Signal_Debounce_0/state[0]_net_1\, 
        \Pressure_Signal_Debounce_0/state[1]_net_1\, 
        Pressure_Signal_Debounce_0_low_pressure, 
        \Science_0/ADC_READ_0/chan[0]_net_1\, 
        \Science_0/ADC_READ_0/chan[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt1dn[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt1dn[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt1dn[2]_net_1\, 
        \Science_0/ADC_READ_0/cnt1dn[3]_net_1\, 
        \Science_0/ADC_READ_0/cnt1dn[4]_net_1\, 
        \Science_0/ADC_READ_0/cnt1dn[5]_net_1\, 
        \Science_0/ADC_READ_0/cnt1dn[6]_net_1\, 
        \Science_0/ADC_READ_0/cnt1dn[7]_net_1\, 
        \Science_0/ADC_READ_0/cnt1up[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt1up[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt1up[2]_net_1\, 
        \Science_0/ADC_READ_0/cnt1up[3]_net_1\, 
        \Science_0/ADC_READ_0/cnt1up[4]_net_1\, 
        \Science_0/ADC_READ_0/cnt2dn[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt2dn[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt2dn[2]_net_1\, 
        \Science_0/ADC_READ_0/cnt2dn[3]_net_1\, 
        \Science_0/ADC_READ_0/cnt2dn[4]_net_1\, 
        \Science_0/ADC_READ_0/cnt2dn[5]_net_1\, 
        \Science_0/ADC_READ_0/cnt2dn[6]_net_1\, 
        \Science_0/ADC_READ_0/cnt2dn[7]_net_1\, 
        \Science_0/ADC_READ_0/cnt2up[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt2up[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt2up[2]_net_1\, 
        \Science_0/ADC_READ_0/cnt2up[3]_net_1\, 
        \Science_0/ADC_READ_0/cnt2up[4]_net_1\, 
        \Science_0/ADC_READ_0/cnt3dn[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt3dn[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt3dn[2]_net_1\, 
        \Science_0/ADC_READ_0/cnt3dn[3]_net_1\, 
        \Science_0/ADC_READ_0/cnt3dn[4]_net_1\, 
        \Science_0/ADC_READ_0/cnt3dn[5]_net_1\, 
        \Science_0/ADC_READ_0/cnt3dn[6]_net_1\, 
        \Science_0/ADC_READ_0/cnt3dn[7]_net_1\, 
        \Science_0/ADC_READ_0/cnt3up[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt3up[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt3up[2]_net_1\, 
        \Science_0/ADC_READ_0/cnt3up[3]_net_1\, 
        \Science_0/ADC_READ_0/cnt3up[4]_net_1\, 
        \Science_0/ADC_READ_0/cnt4dn[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt4dn[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt4dn[2]_net_1\, 
        \Science_0/ADC_READ_0/cnt4dn[3]_net_1\, 
        \Science_0/ADC_READ_0/cnt4dn[4]_net_1\, 
        \Science_0/ADC_READ_0/cnt4dn[5]_net_1\, 
        \Science_0/ADC_READ_0/cnt4dn[6]_net_1\, 
        \Science_0/ADC_READ_0/cnt4dn[7]_net_1\, 
        \Science_0/ADC_READ_0/cnt4up[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt4up[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt4up[2]_net_1\, 
        \Science_0/ADC_READ_0/cnt4up[3]_net_1\, 
        \Science_0/ADC_READ_0/cnt4up[4]_net_1\, 
        \Science_0/ADC_READ_0/cnt[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt[1]_net_1\, 
        \Science_0/ADC_READ_0/cnt[2]_net_1\, 
        \Science_0/ADC_READ_0/cnt[3]_net_1\, 
        \Science_0/ADC_READ_0/cnt[4]_net_1\, 
        \Science_0/ADC_READ_0/cnt[5]_net_1\, 
        \Science_0/ADC_READ_0/cnt[6]_net_1\, 
        \Science_0/ADC_READ_0/cnt[7]_net_1\, 
        \Science_0/ADC_READ_0/cnt_chan[0]_net_1\, 
        \Science_0/ADC_READ_0/cnt_chan[1]_net_1\, 
        \Science_0/ADC_READ_0/countere\, 
        \Science_0/ADC_READ_0/data_a[0]_net_1\, 
        \Science_0/ADC_READ_0/data_a[10]_net_1\, 
        \Science_0/ADC_READ_0/data_a[11]_net_1\, 
        \Science_0/ADC_READ_0/data_a[12]_net_1\, 
        \Science_0/ADC_READ_0/data_a[13]_net_1\, 
        \Science_0/ADC_READ_0/data_a[14]_net_1\, 
        \Science_0/ADC_READ_0/data_a[15]_net_1\, 
        \Science_0/ADC_READ_0/data_a[16]_net_1\, 
        \Science_0/ADC_READ_0/data_a[17]_net_1\, 
        \Science_0/ADC_READ_0/data_a[1]_net_1\, 
        \Science_0/ADC_READ_0/data_a[2]_net_1\, 
        \Science_0/ADC_READ_0/data_a[3]_net_1\, 
        \Science_0/ADC_READ_0/data_a[4]_net_1\, 
        \Science_0/ADC_READ_0/data_a[5]_net_1\, 
        \Science_0/ADC_READ_0/data_a[6]_net_1\, 
        \Science_0/ADC_READ_0/data_a[7]_net_1\, 
        \Science_0/ADC_READ_0/data_a[8]_net_1\, 
        \Science_0/ADC_READ_0/data_a[9]_net_1\, 
        \Science_0/ADC_READ_0/data_b[0]_net_1\, 
        \Science_0/ADC_READ_0/data_b[10]_net_1\, 
        \Science_0/ADC_READ_0/data_b[11]_net_1\, 
        \Science_0/ADC_READ_0/data_b[12]_net_1\, 
        \Science_0/ADC_READ_0/data_b[13]_net_1\, 
        \Science_0/ADC_READ_0/data_b[14]_net_1\, 
        \Science_0/ADC_READ_0/data_b[15]_net_1\, 
        \Science_0/ADC_READ_0/data_b[16]_net_1\, 
        \Science_0/ADC_READ_0/data_b[17]_net_1\, 
        \Science_0/ADC_READ_0/data_b[1]_net_1\, 
        \Science_0/ADC_READ_0/data_b[2]_net_1\, 
        \Science_0/ADC_READ_0/data_b[3]_net_1\, 
        \Science_0/ADC_READ_0/data_b[4]_net_1\, 
        \Science_0/ADC_READ_0/data_b[5]_net_1\, 
        \Science_0/ADC_READ_0/data_b[6]_net_1\, 
        \Science_0/ADC_READ_0/data_b[7]_net_1\, 
        \Science_0/ADC_READ_0/data_b[8]_net_1\, 
        \Science_0/ADC_READ_0/data_b[9]_net_1\, 
        \Science_0/ADC_READ_0/newflag_net_1\, 
        \Science_0/ADC_READ_0/state[0]_net_1\, 
        \Science_0/ADC_READ_0/state[1]_net_1\, 
        \Science_0/ADC_READ_0/state[2]_net_1\, 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, 
        \Science_0/ADC_READ_0_G1[0]\, 
        \Science_0/ADC_READ_0_G1[1]\, 
        \Science_0/ADC_READ_0_G2[0]\, 
        \Science_0/ADC_READ_0_G2[1]\, 
        \Science_0/ADC_READ_0_G3[0]\, 
        \Science_0/ADC_READ_0_G3[1]\, 
        \Science_0/ADC_READ_0_G4[0]\, 
        \Science_0/ADC_READ_0_G4[1]\, 
        \Science_0/ADC_RESET_0/old_enable_net_1\, 
        \Science_0/ADC_RESET_0/state[0]_net_1\, 
        \Science_0/ADC_RESET_0/state[1]_net_1\, 
        \Science_0/DAC_SET_0/ADR[0]_net_1\, 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, 
        \Science_0/DAC_SET_0/cnt[0]_net_1\, 
        \Science_0/DAC_SET_0/cnt[1]_net_1\, 
        \Science_0/DAC_SET_0/cnt[2]_net_1\, 
        \Science_0/DAC_SET_0/cnt[3]_net_1\, 
        \Science_0/DAC_SET_0/cnt[4]_net_1\, 
        \Science_0/DAC_SET_0/old_set_net_1\, 
        \Science_0/DAC_SET_0/state[1]_net_1\, 
        \Science_0/DAC_SET_0/state[2]_net_1\, 
        \Science_0/DAC_SET_0/state[3]_net_1\, 
        \Science_0/DAC_SET_0/state[4]_net_1\, 
        \Science_0/DAC_SET_0/vector[0]_net_1\, 
        \Science_0/DAC_SET_0/vector[10]_net_1\, 
        \Science_0/DAC_SET_0/vector[11]_net_1\, 
        \Science_0/DAC_SET_0/vector[12]_net_1\, 
        \Science_0/DAC_SET_0/vector[13]_net_1\, 
        \Science_0/DAC_SET_0/vector[14]_net_1\, 
        \Science_0/DAC_SET_0/vector[15]_net_1\, 
        \Science_0/DAC_SET_0/vector[16]_net_1\, 
        \Science_0/DAC_SET_0/vector[17]_net_1\, 
        \Science_0/DAC_SET_0/vector[1]_net_1\, 
        \Science_0/DAC_SET_0/vector[2]_net_1\, 
        \Science_0/DAC_SET_0/vector[3]_net_1\, 
        \Science_0/DAC_SET_0/vector[4]_net_1\, 
        \Science_0/DAC_SET_0/vector[5]_net_1\, 
        \Science_0/DAC_SET_0/vector[6]_net_1\, 
        \Science_0/DAC_SET_0/vector[7]_net_1\, 
        \Science_0/DAC_SET_0/vector[8]_net_1\, 
        \Science_0/DAC_SET_0/vector[9]_net_1\, 
        \Science_0/SET_LP_GAIN_0/old_G1[0]_net_1\, 
        \Science_0/SET_LP_GAIN_0/old_G1[1]_net_1\, 
        \Science_0/SET_LP_GAIN_0/old_G2[0]_net_1\, 
        \Science_0/SET_LP_GAIN_0/old_G2[1]_net_1\, 
        \Science_0/SET_LP_GAIN_0/old_G3[0]_net_1\, 
        \Science_0/SET_LP_GAIN_0/old_G3[1]_net_1\, 
        \Science_0/SET_LP_GAIN_0/old_G4[0]_net_1\, 
        \Science_0/SET_LP_GAIN_0/old_G4[1]_net_1\, 
        \Science_0/SET_LP_GAIN_0/state[4]_net_1\, 
        \Science_0/SET_LP_GAIN_0/state[5]_net_1\, 
        \Science_0/SET_LP_GAIN_0/state[6]_net_1\, 
        \Science_0/SET_LP_GAIN_0/state[7]_net_1\, 
        \Science_0/SET_LP_GAIN_0/state_i_0[0]\, 
        \Science_0/SET_LP_GAIN_0/state_i_0[1]\, 
        \Science_0/SET_LP_GAIN_0/state_i_0[2]\, 
        \Science_0/SET_LP_GAIN_0/state_i_0[3]\, 
        \Science_0/SWEEP_SPIDER2_0/latch_i_0\, 
        \Science_0/SWEEP_SPIDER2_0_SET\, 
        \Science_0_chan0_data[0]\, \Science_0_chan0_data[10]\, 
        \Science_0_chan0_data[11]\, \Science_0_chan0_data[1]\, 
        \Science_0_chan0_data[2]\, \Science_0_chan0_data[3]\, 
        \Science_0_chan0_data[4]\, \Science_0_chan0_data[5]\, 
        \Science_0_chan0_data[6]\, \Science_0_chan0_data[7]\, 
        \Science_0_chan0_data[8]\, \Science_0_chan0_data[9]\, 
        \Science_0_chan1_data[0]\, \Science_0_chan1_data[10]\, 
        \Science_0_chan1_data[11]\, \Science_0_chan1_data[1]\, 
        \Science_0_chan1_data[2]\, \Science_0_chan1_data[3]\, 
        \Science_0_chan1_data[4]\, \Science_0_chan1_data[5]\, 
        \Science_0_chan1_data[6]\, \Science_0_chan1_data[7]\, 
        \Science_0_chan1_data[8]\, \Science_0_chan1_data[9]\, 
        \Science_0_chan2_data[0]\, \Science_0_chan2_data[10]\, 
        \Science_0_chan2_data[11]\, \Science_0_chan2_data[1]\, 
        \Science_0_chan2_data[2]\, \Science_0_chan2_data[3]\, 
        \Science_0_chan2_data[4]\, \Science_0_chan2_data[5]\, 
        \Science_0_chan2_data[6]\, \Science_0_chan2_data[7]\, 
        \Science_0_chan2_data[8]\, \Science_0_chan2_data[9]\, 
        \Science_0_chan3_data[0]\, \Science_0_chan3_data[10]\, 
        \Science_0_chan3_data[11]\, \Science_0_chan3_data[1]\, 
        \Science_0_chan3_data[2]\, \Science_0_chan3_data[3]\, 
        \Science_0_chan3_data[4]\, \Science_0_chan3_data[5]\, 
        \Science_0_chan3_data[6]\, \Science_0_chan3_data[7]\, 
        \Science_0_chan3_data[8]\, \Science_0_chan3_data[9]\, 
        \Science_0_chan4_data[0]\, \Science_0_chan4_data[10]\, 
        \Science_0_chan4_data[11]\, \Science_0_chan4_data[1]\, 
        \Science_0_chan4_data[2]\, \Science_0_chan4_data[3]\, 
        \Science_0_chan4_data[4]\, \Science_0_chan4_data[5]\, 
        \Science_0_chan4_data[6]\, \Science_0_chan4_data[7]\, 
        \Science_0_chan4_data[8]\, \Science_0_chan4_data[9]\, 
        \Science_0_chan5_data[0]\, \Science_0_chan5_data[10]\, 
        \Science_0_chan5_data[11]\, \Science_0_chan5_data[1]\, 
        \Science_0_chan5_data[2]\, \Science_0_chan5_data[3]\, 
        \Science_0_chan5_data[4]\, \Science_0_chan5_data[5]\, 
        \Science_0_chan5_data[6]\, \Science_0_chan5_data[7]\, 
        \Science_0_chan5_data[8]\, \Science_0_chan5_data[9]\, 
        \Science_0_chan6_data[0]\, \Science_0_chan6_data[10]\, 
        \Science_0_chan6_data[11]\, \Science_0_chan6_data[1]\, 
        \Science_0_chan6_data[2]\, \Science_0_chan6_data[3]\, 
        \Science_0_chan6_data[4]\, \Science_0_chan6_data[5]\, 
        \Science_0_chan6_data[6]\, \Science_0_chan6_data[7]\, 
        \Science_0_chan6_data[8]\, \Science_0_chan6_data[9]\, 
        \Science_0_chan7_data[0]\, \Science_0_chan7_data[10]\, 
        \Science_0_chan7_data[11]\, \Science_0_chan7_data[1]\, 
        \Science_0_chan7_data[2]\, \Science_0_chan7_data[3]\, 
        \Science_0_chan7_data[4]\, \Science_0_chan7_data[5]\, 
        \Science_0_chan7_data[6]\, \Science_0_chan7_data[7]\, 
        \Science_0_chan7_data[8]\, \Science_0_chan7_data[9]\, 
        Science_0_exp_new_data, \Science_0_exp_packet_0[0]\, 
        \Science_0_exp_packet_0[11]\, 
        \Science_0_exp_packet_0[12]\, 
        \Science_0_exp_packet_0[15]\, 
        \Science_0_exp_packet_0[16]\, 
        \Science_0_exp_packet_0[17]\, 
        \Science_0_exp_packet_0[18]\, 
        \Science_0_exp_packet_0[19]\, \Science_0_exp_packet_0[1]\, 
        \Science_0_exp_packet_0[20]\, 
        \Science_0_exp_packet_0[21]\, 
        \Science_0_exp_packet_0[22]\, 
        \Science_0_exp_packet_0[23]\, 
        \Science_0_exp_packet_0[24]\, 
        \Science_0_exp_packet_0[25]\, 
        \Science_0_exp_packet_0[26]\, 
        \Science_0_exp_packet_0[27]\, 
        \Science_0_exp_packet_0[28]\, 
        \Science_0_exp_packet_0[29]\, \Science_0_exp_packet_0[2]\, 
        \Science_0_exp_packet_0[30]\, 
        \Science_0_exp_packet_0[31]\, 
        \Science_0_exp_packet_0[32]\, 
        \Science_0_exp_packet_0[33]\, 
        \Science_0_exp_packet_0[34]\, 
        \Science_0_exp_packet_0[35]\, 
        \Science_0_exp_packet_0[36]\, 
        \Science_0_exp_packet_0[37]\, 
        \Science_0_exp_packet_0[38]\, 
        \Science_0_exp_packet_0[39]\, \Science_0_exp_packet_0[3]\, 
        \Science_0_exp_packet_0[40]\, 
        \Science_0_exp_packet_0[41]\, 
        \Science_0_exp_packet_0[42]\, 
        \Science_0_exp_packet_0[43]\, 
        \Science_0_exp_packet_0[44]\, 
        \Science_0_exp_packet_0[45]\, 
        \Science_0_exp_packet_0[46]\, 
        \Science_0_exp_packet_0[47]\, 
        \Science_0_exp_packet_0[48]\, 
        \Science_0_exp_packet_0[49]\, \Science_0_exp_packet_0[4]\, 
        \Science_0_exp_packet_0[50]\, 
        \Science_0_exp_packet_0[51]\, 
        \Science_0_exp_packet_0[52]\, 
        \Science_0_exp_packet_0[53]\, 
        \Science_0_exp_packet_0[54]\, 
        \Science_0_exp_packet_0[55]\, 
        \Science_0_exp_packet_0[56]\, 
        \Science_0_exp_packet_0[57]\, 
        \Science_0_exp_packet_0[58]\, 
        \Science_0_exp_packet_0[59]\, 
        \Science_0_exp_packet_0[60]\, 
        \Science_0_exp_packet_0[61]\, 
        \Science_0_exp_packet_0[62]\, 
        \Science_0_exp_packet_0[63]\, 
        \Science_0_exp_packet_0[64]\, 
        \Science_0_exp_packet_0[65]\, 
        \Science_0_exp_packet_0[66]\, 
        \Science_0_exp_packet_0[67]\, 
        \Science_0_exp_packet_0[68]\, 
        \Science_0_exp_packet_0[69]\, 
        \Science_0_exp_packet_0[70]\, 
        \Science_0_exp_packet_0[71]\, 
        \Science_0_exp_packet_0[72]\, 
        \Science_0_exp_packet_0[73]\, 
        \Science_0_exp_packet_0[74]\, 
        \Science_0_exp_packet_0[75]\, 
        \Science_0_exp_packet_0[76]\, 
        \Science_0_exp_packet_0[77]\, 
        \Science_0_exp_packet_0[78]\, 
        \Science_0_exp_packet_0[79]\, \Science_0_exp_packet_0[8]\, 
        \Science_0_exp_packet_0[9]\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[3]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[2]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[3]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_1_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_2_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/isSetup_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[0]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[1]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[2]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[3]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[4]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[5]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[6]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[7]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[8]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[3]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[0]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[2]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[3]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[4]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[5]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[6]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[7]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[0]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[1]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[2]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[3]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_repeat_start\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[0]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[1]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[2]\, 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_we\, 
        \Sensors_0/Accelerometer_0/state[8]\, 
        \Sensors_0/Accelerometer_0/state_0[8]\, 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[2]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[3]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[0]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_1_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_2_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/state[2]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/state[5]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[0]\, 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[1]\, 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[2]\, 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[4]\, 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[5]\, 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[6]\, 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[7]\, 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, 
        \Sensors_0/Gyro_0/I2C_Master_0_s_ack_error\, 
        \Sensors_0/Gyro_0/I2C_Master_0_write_done\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/isSetup_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[1]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[2]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[3]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[5]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[6]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[7]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[0]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[1]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[2]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[3]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[6]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[7]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_i2c_addr[0]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_i2c_repeat_start\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_num_bytes[0]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_num_bytes[1]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_num_bytes[2]\, 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_we\, 
        \Sensors_0/Gyro_0/state[8]\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[2]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[3]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[0]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[2]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_1_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_2_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[2]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[5]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[0]\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[1]\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[2]\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[3]\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[4]\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[5]\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[6]\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[7]\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_s_ack_error\, 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_write_done\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/isSetup_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[0]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[1]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[2]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[3]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[4]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[5]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[6]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[7]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[1]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[3]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[2]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[4]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[5]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[1]\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[3]\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[4]\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[6]\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_i2c_addr[0]\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_num_bytes[0]\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_num_bytes[1]\, 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_we\, 
        \Sensors_0/Pressure_Sensor_0/state[8]\, 
        Sensors_0_acc_new_data, \Sensors_0_acc_temp[0]\, 
        \Sensors_0_acc_temp[1]\, \Sensors_0_acc_temp[2]\, 
        \Sensors_0_acc_temp[3]\, \Sensors_0_acc_temp[4]\, 
        \Sensors_0_acc_temp[5]\, \Sensors_0_acc_temp[6]\, 
        \Sensors_0_acc_temp[7]\, \Sensors_0_acc_time[0]\, 
        \Sensors_0_acc_time[10]\, \Sensors_0_acc_time[11]\, 
        \Sensors_0_acc_time[12]\, \Sensors_0_acc_time[13]\, 
        \Sensors_0_acc_time[14]\, \Sensors_0_acc_time[15]\, 
        \Sensors_0_acc_time[16]\, \Sensors_0_acc_time[17]\, 
        \Sensors_0_acc_time[18]\, \Sensors_0_acc_time[19]\, 
        \Sensors_0_acc_time[1]\, \Sensors_0_acc_time[20]\, 
        \Sensors_0_acc_time[21]\, \Sensors_0_acc_time[22]\, 
        \Sensors_0_acc_time[23]\, \Sensors_0_acc_time[2]\, 
        \Sensors_0_acc_time[3]\, \Sensors_0_acc_time[4]\, 
        \Sensors_0_acc_time[5]\, \Sensors_0_acc_time[6]\, 
        \Sensors_0_acc_time[7]\, \Sensors_0_acc_time[8]\, 
        \Sensors_0_acc_time[9]\, \Sensors_0_acc_x[0]\, 
        \Sensors_0_acc_x[10]\, \Sensors_0_acc_x[11]\, 
        \Sensors_0_acc_x[1]\, \Sensors_0_acc_x[2]\, 
        \Sensors_0_acc_x[3]\, \Sensors_0_acc_x[4]\, 
        \Sensors_0_acc_x[5]\, \Sensors_0_acc_x[6]\, 
        \Sensors_0_acc_x[7]\, \Sensors_0_acc_x[8]\, 
        \Sensors_0_acc_x[9]\, \Sensors_0_acc_y[0]\, 
        \Sensors_0_acc_y[10]\, \Sensors_0_acc_y[11]\, 
        \Sensors_0_acc_y[1]\, \Sensors_0_acc_y[2]\, 
        \Sensors_0_acc_y[3]\, \Sensors_0_acc_y[4]\, 
        \Sensors_0_acc_y[5]\, \Sensors_0_acc_y[6]\, 
        \Sensors_0_acc_y[7]\, \Sensors_0_acc_y[8]\, 
        \Sensors_0_acc_y[9]\, \Sensors_0_acc_z[0]\, 
        \Sensors_0_acc_z[10]\, \Sensors_0_acc_z[11]\, 
        \Sensors_0_acc_z[1]\, \Sensors_0_acc_z[2]\, 
        \Sensors_0_acc_z[3]\, \Sensors_0_acc_z[4]\, 
        \Sensors_0_acc_z[5]\, \Sensors_0_acc_z[6]\, 
        \Sensors_0_acc_z[7]\, \Sensors_0_acc_z[8]\, 
        \Sensors_0_acc_z[9]\, Sensors_0_gyro_new_data, 
        \Sensors_0_gyro_temp[0]\, \Sensors_0_gyro_temp[1]\, 
        \Sensors_0_gyro_temp[2]\, \Sensors_0_gyro_temp[3]\, 
        \Sensors_0_gyro_temp[4]\, \Sensors_0_gyro_temp[5]\, 
        \Sensors_0_gyro_temp[6]\, \Sensors_0_gyro_temp[7]\, 
        \Sensors_0_gyro_time[0]\, \Sensors_0_gyro_time[10]\, 
        \Sensors_0_gyro_time[11]\, \Sensors_0_gyro_time[12]\, 
        \Sensors_0_gyro_time[13]\, \Sensors_0_gyro_time[14]\, 
        \Sensors_0_gyro_time[15]\, \Sensors_0_gyro_time[16]\, 
        \Sensors_0_gyro_time[17]\, \Sensors_0_gyro_time[18]\, 
        \Sensors_0_gyro_time[19]\, \Sensors_0_gyro_time[1]\, 
        \Sensors_0_gyro_time[20]\, \Sensors_0_gyro_time[21]\, 
        \Sensors_0_gyro_time[22]\, \Sensors_0_gyro_time[23]\, 
        \Sensors_0_gyro_time[2]\, \Sensors_0_gyro_time[3]\, 
        \Sensors_0_gyro_time[4]\, \Sensors_0_gyro_time[5]\, 
        \Sensors_0_gyro_time[6]\, \Sensors_0_gyro_time[7]\, 
        \Sensors_0_gyro_time[8]\, \Sensors_0_gyro_time[9]\, 
        \Sensors_0_gyro_x[0]\, \Sensors_0_gyro_x[10]\, 
        \Sensors_0_gyro_x[11]\, \Sensors_0_gyro_x[12]\, 
        \Sensors_0_gyro_x[13]\, \Sensors_0_gyro_x[14]\, 
        \Sensors_0_gyro_x[15]\, \Sensors_0_gyro_x[1]\, 
        \Sensors_0_gyro_x[2]\, \Sensors_0_gyro_x[3]\, 
        \Sensors_0_gyro_x[4]\, \Sensors_0_gyro_x[5]\, 
        \Sensors_0_gyro_x[6]\, \Sensors_0_gyro_x[7]\, 
        \Sensors_0_gyro_x[8]\, \Sensors_0_gyro_x[9]\, 
        \Sensors_0_gyro_y[0]\, \Sensors_0_gyro_y[10]\, 
        \Sensors_0_gyro_y[11]\, \Sensors_0_gyro_y[12]\, 
        \Sensors_0_gyro_y[13]\, \Sensors_0_gyro_y[14]\, 
        \Sensors_0_gyro_y[15]\, \Sensors_0_gyro_y[1]\, 
        \Sensors_0_gyro_y[2]\, \Sensors_0_gyro_y[3]\, 
        \Sensors_0_gyro_y[4]\, \Sensors_0_gyro_y[5]\, 
        \Sensors_0_gyro_y[6]\, \Sensors_0_gyro_y[7]\, 
        \Sensors_0_gyro_y[8]\, \Sensors_0_gyro_y[9]\, 
        \Sensors_0_gyro_z[0]\, \Sensors_0_gyro_z[1]\, 
        \Sensors_0_gyro_z[2]\, \Sensors_0_gyro_z[3]\, 
        Sensors_0_mag_new_data, \Sensors_0_mag_time[0]\, 
        \Sensors_0_mag_time[10]\, \Sensors_0_mag_time[11]\, 
        \Sensors_0_mag_time[12]\, \Sensors_0_mag_time[13]\, 
        \Sensors_0_mag_time[14]\, \Sensors_0_mag_time[15]\, 
        \Sensors_0_mag_time[16]\, \Sensors_0_mag_time[17]\, 
        \Sensors_0_mag_time[18]\, \Sensors_0_mag_time[19]\, 
        \Sensors_0_mag_time[1]\, \Sensors_0_mag_time[20]\, 
        \Sensors_0_mag_time[21]\, \Sensors_0_mag_time[22]\, 
        \Sensors_0_mag_time[23]\, \Sensors_0_mag_time[2]\, 
        \Sensors_0_mag_time[3]\, \Sensors_0_mag_time[4]\, 
        \Sensors_0_mag_time[5]\, \Sensors_0_mag_time[6]\, 
        \Sensors_0_mag_time[7]\, \Sensors_0_mag_time[8]\, 
        \Sensors_0_mag_time[9]\, \Sensors_0_mag_x[0]\, 
        \Sensors_0_mag_x[10]\, \Sensors_0_mag_x[11]\, 
        \Sensors_0_mag_x[1]\, \Sensors_0_mag_x[2]\, 
        \Sensors_0_mag_x[3]\, \Sensors_0_mag_x[4]\, 
        \Sensors_0_mag_x[5]\, \Sensors_0_mag_x[6]\, 
        \Sensors_0_mag_x[7]\, \Sensors_0_mag_x[8]\, 
        \Sensors_0_mag_x[9]\, \Sensors_0_mag_y[0]\, 
        \Sensors_0_mag_y[10]\, \Sensors_0_mag_y[11]\, 
        \Sensors_0_mag_y[1]\, \Sensors_0_mag_y[2]\, 
        \Sensors_0_mag_y[3]\, \Sensors_0_mag_y[4]\, 
        \Sensors_0_mag_y[5]\, \Sensors_0_mag_y[6]\, 
        \Sensors_0_mag_y[7]\, \Sensors_0_mag_y[8]\, 
        \Sensors_0_mag_y[9]\, \Sensors_0_mag_z[0]\, 
        \Sensors_0_mag_z[10]\, \Sensors_0_mag_z[11]\, 
        \Sensors_0_mag_z[1]\, \Sensors_0_mag_z[2]\, 
        \Sensors_0_mag_z[3]\, \Sensors_0_mag_z[4]\, 
        \Sensors_0_mag_z[5]\, \Sensors_0_mag_z[6]\, 
        \Sensors_0_mag_z[7]\, \Sensors_0_mag_z[8]\, 
        \Sensors_0_mag_z[9]\, Sensors_0_pressure_new_data, 
        \Sensors_0_pressure_raw[0]\, \Sensors_0_pressure_raw[10]\, 
        \Sensors_0_pressure_raw[11]\, 
        \Sensors_0_pressure_raw[12]\, 
        \Sensors_0_pressure_raw[13]\, 
        \Sensors_0_pressure_raw[14]\, 
        \Sensors_0_pressure_raw[15]\, 
        \Sensors_0_pressure_raw[16]\, 
        \Sensors_0_pressure_raw[17]\, 
        \Sensors_0_pressure_raw[18]\, 
        \Sensors_0_pressure_raw[19]\, \Sensors_0_pressure_raw[1]\, 
        \Sensors_0_pressure_raw[20]\, 
        \Sensors_0_pressure_raw[21]\, 
        \Sensors_0_pressure_raw[22]\, 
        \Sensors_0_pressure_raw[23]\, \Sensors_0_pressure_raw[2]\, 
        \Sensors_0_pressure_raw[3]\, \Sensors_0_pressure_raw[4]\, 
        \Sensors_0_pressure_raw[5]\, \Sensors_0_pressure_raw[6]\, 
        \Sensors_0_pressure_raw[7]\, \Sensors_0_pressure_raw[8]\, 
        \Sensors_0_pressure_raw[9]\, 
        \Sensors_0_pressure_temp_raw[0]\, 
        \Sensors_0_pressure_temp_raw[10]\, 
        \Sensors_0_pressure_temp_raw[11]\, 
        \Sensors_0_pressure_temp_raw[12]\, 
        \Sensors_0_pressure_temp_raw[13]\, 
        \Sensors_0_pressure_temp_raw[14]\, 
        \Sensors_0_pressure_temp_raw[15]\, 
        \Sensors_0_pressure_temp_raw[16]\, 
        \Sensors_0_pressure_temp_raw[17]\, 
        \Sensors_0_pressure_temp_raw[18]\, 
        \Sensors_0_pressure_temp_raw[19]\, 
        \Sensors_0_pressure_temp_raw[1]\, 
        \Sensors_0_pressure_temp_raw[20]\, 
        \Sensors_0_pressure_temp_raw[21]\, 
        \Sensors_0_pressure_temp_raw[22]\, 
        \Sensors_0_pressure_temp_raw[23]\, 
        \Sensors_0_pressure_temp_raw[2]\, 
        \Sensors_0_pressure_temp_raw[3]\, 
        \Sensors_0_pressure_temp_raw[4]\, 
        \Sensors_0_pressure_temp_raw[5]\, 
        \Sensors_0_pressure_temp_raw[6]\, 
        \Sensors_0_pressure_temp_raw[7]\, 
        \Sensors_0_pressure_temp_raw[8]\, 
        \Sensors_0_pressure_temp_raw[9]\, 
        \Sensors_0_pressure_time[0]\, 
        \Sensors_0_pressure_time[10]\, 
        \Sensors_0_pressure_time[11]\, 
        \Sensors_0_pressure_time[12]\, 
        \Sensors_0_pressure_time[13]\, 
        \Sensors_0_pressure_time[14]\, 
        \Sensors_0_pressure_time[15]\, 
        \Sensors_0_pressure_time[16]\, 
        \Sensors_0_pressure_time[17]\, 
        \Sensors_0_pressure_time[18]\, 
        \Sensors_0_pressure_time[19]\, 
        \Sensors_0_pressure_time[1]\, 
        \Sensors_0_pressure_time[20]\, 
        \Sensors_0_pressure_time[21]\, 
        \Sensors_0_pressure_time[22]\, 
        \Sensors_0_pressure_time[23]\, 
        \Sensors_0_pressure_time[2]\, 
        \Sensors_0_pressure_time[3]\, 
        \Sensors_0_pressure_time[4]\, 
        \Sensors_0_pressure_time[5]\, 
        \Sensors_0_pressure_time[6]\, 
        \Sensors_0_pressure_time[7]\, 
        \Sensors_0_pressure_time[8]\, 
        \Sensors_0_pressure_time[9]\, 
        \Timekeeper_0/old_1MHz_net_1\, 
        \Timekeeper_0/old_1kHz_net_1\, 
        \Timekeeper_0_microseconds[0]\, 
        \Timekeeper_0_microseconds[10]\, 
        \Timekeeper_0_microseconds[11]\, 
        \Timekeeper_0_microseconds[12]\, 
        \Timekeeper_0_microseconds[13]\, 
        \Timekeeper_0_microseconds[14]\, 
        \Timekeeper_0_microseconds[15]\, 
        \Timekeeper_0_microseconds[16]\, 
        \Timekeeper_0_microseconds[17]\, 
        \Timekeeper_0_microseconds[18]\, 
        \Timekeeper_0_microseconds[19]\, 
        \Timekeeper_0_microseconds[1]\, 
        \Timekeeper_0_microseconds[20]\, 
        \Timekeeper_0_microseconds[21]\, 
        \Timekeeper_0_microseconds[22]\, 
        \Timekeeper_0_microseconds[23]\, 
        \Timekeeper_0_microseconds[2]\, 
        \Timekeeper_0_microseconds[3]\, 
        \Timekeeper_0_microseconds[4]\, 
        \Timekeeper_0_microseconds[5]\, 
        \Timekeeper_0_microseconds[6]\, 
        \Timekeeper_0_microseconds[7]\, 
        \Timekeeper_0_microseconds[8]\, 
        \Timekeeper_0_microseconds[9]\, 
        \Timekeeper_0_milliseconds[0]\, 
        \Timekeeper_0_milliseconds[10]\, 
        \Timekeeper_0_milliseconds[11]\, 
        \Timekeeper_0_milliseconds[12]\, 
        \Timekeeper_0_milliseconds[13]\, 
        \Timekeeper_0_milliseconds[14]\, 
        \Timekeeper_0_milliseconds[15]\, 
        \Timekeeper_0_milliseconds[16]\, 
        \Timekeeper_0_milliseconds[17]\, 
        \Timekeeper_0_milliseconds[18]\, 
        \Timekeeper_0_milliseconds[19]\, 
        \Timekeeper_0_milliseconds[1]\, 
        \Timekeeper_0_milliseconds[20]\, 
        \Timekeeper_0_milliseconds[21]\, 
        \Timekeeper_0_milliseconds[22]\, 
        \Timekeeper_0_milliseconds[23]\, 
        \Timekeeper_0_milliseconds[2]\, 
        \Timekeeper_0_milliseconds[3]\, 
        \Timekeeper_0_milliseconds[4]\, 
        \Timekeeper_0_milliseconds[5]\, 
        \Timekeeper_0_milliseconds[6]\, 
        \Timekeeper_0_milliseconds[7]\, 
        \Timekeeper_0_milliseconds[8]\, 
        \Timekeeper_0_milliseconds[9]\, 
        \Timing_0/f_time[0]_net_1\, \Timing_0/f_time[1]_net_1\, 
        \Timing_0/f_time[2]_net_1\, \Timing_0/f_time[3]_net_1\, 
        \Timing_0/m_count[0]_net_1\, \Timing_0/m_count[1]_net_1\, 
        \Timing_0/m_count[2]_net_1\, \Timing_0/m_count[3]_net_1\, 
        \Timing_0/m_count[4]_net_1\, \Timing_0/m_count[5]_net_1\, 
        \Timing_0/m_count[6]_net_1\, \Timing_0/m_count[7]_net_1\, 
        \Timing_0/m_time[0]_net_1\, \Timing_0/m_time[1]_net_1\, 
        \Timing_0/m_time[3]_net_1\, \Timing_0/m_time[4]_net_1\, 
        \Timing_0/m_time[5]_net_1\, \Timing_0/m_time[6]_net_1\, 
        \Timing_0/s_count[0]_net_1\, \Timing_0/s_count[1]_net_1\, 
        \Timing_0/s_count[2]_net_1\, \Timing_0/s_count[3]_net_1\, 
        \Timing_0/s_count[4]_net_1\, \Timing_0/s_count[5]_net_1\, 
        \Timing_0/s_count[6]_net_1\, \Timing_0/s_count[7]_net_1\, 
        \Timing_0/s_time[0]_net_1\, \Timing_0/s_time[1]_net_1\, 
        \Timing_0/s_time[2]_net_1\, \Timing_0/s_time[4]_net_1\, 
        \Timing_0/s_time[6]_net_1\, \Timing_0/s_time[7]_net_1\, 
        \Timing_0/s_time[8]_net_1\, \ch3_data_net_0[0]\, 
        \ch3_data_net_0[10]\, \ch3_data_net_0[11]\, 
        \ch3_data_net_0[1]\, \ch3_data_net_0[2]\, 
        \ch3_data_net_0[3]\, \ch3_data_net_0[4]\, 
        \ch3_data_net_0[5]\, \ch3_data_net_0[6]\, 
        \ch3_data_net_0[7]\, \ch3_data_net_0[8]\, 
        \ch3_data_net_0[9]\, \m_time[7]\, \s_clks_net_0[18]\, 
        \s_clks_net_0[24]\, \s_clks_net_0[4]\, \s_clks_net_0[9]\, 
        \s_time[5]\, AFLSDF_VCC, AFLSDF_GND, \AFLSDF_INV_0\, 
        \AFLSDF_INV_1\, \AFLSDF_INV_2\, \AFLSDF_INV_3\, 
        \AFLSDF_INV_4\, \AFLSDF_INV_5\, \AFLSDF_INV_6\, 
        \AFLSDF_INV_7\, \AFLSDF_INV_8\, \AFLSDF_INV_9\, 
        \AFLSDF_INV_10\, \AFLSDF_INV_11\, \AFLSDF_INV_12\, 
        \AFLSDF_INV_13\, \AFLSDF_INV_14\, \AFLSDF_INV_15\, 
        \AFLSDF_INV_16\, \AFLSDF_INV_17\, \AFLSDF_INV_18\, 
        \AFLSDF_INV_19\, \AFLSDF_INV_20\, \AFLSDF_INV_21\, 
        \AFLSDF_INV_22\, \AFLSDF_INV_23\, \AFLSDF_INV_24\, 
        \AFLSDF_INV_25\, \AFLSDF_INV_26\, \AFLSDF_INV_27\, 
        \AFLSDF_INV_28\, \AFLSDF_INV_29\, \AFLSDF_INV_30\, 
        \AFLSDF_INV_31\, \AFLSDF_INV_32\, \AFLSDF_INV_33\, 
        \AFLSDF_INV_34\, \AFLSDF_INV_35\, \AFLSDF_INV_36\, 
        \AFLSDF_INV_37\ : std_logic;
    signal GND_power_net1 : std_logic;
    signal VCC_power_net1 : std_logic;

begin 

    AFLSDF_GND <= GND_power_net1;
    \GND\ <= GND_power_net1;
    \VCC\ <= VCC_power_net1;
    AFLSDF_VCC <= VCC_power_net1;

    \GS_Readout_0/send[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74708, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74630, Q => 
        \GS_Readout_0_send[7]\);
    
    HIEFFPLA_INST_0_61841 : OR3B
      port map(A => HIEFFPLA_NET_0_74117, B => 
        HIEFFPLA_NET_0_74107, C => HIEFFPLA_NET_0_74116, Y => 
        HIEFFPLA_NET_0_74118);
    
    HIEFFPLA_INST_0_66792 : AO1A
      port map(A => HIEFFPLA_NET_0_73098, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73034);
    
    \Data_Saving_0/Packet_Saver_0/data_out[15]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75230, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[15]\);
    
    HIEFFPLA_INST_0_55645 : XA1
      port map(A => \Communications_0/UART_1/rx_clk_count_c0\, B
         => \Communications_0/UART_1/rx_clk_count[30]_net_1\, C
         => HIEFFPLA_NET_0_75437, Y => HIEFFPLA_NET_0_75457);
    
    HIEFFPLA_INST_0_69711 : AOI1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_72322, C => PRESSURE_SCL_c, Y => 
        HIEFFPLA_NET_0_72323);
    
    HIEFFPLA_INST_0_59051 : AO1B
      port map(A => HIEFFPLA_NET_0_74622, B => 
        HIEFFPLA_NET_0_74627, C => HIEFFPLA_NET_0_74625, Y => 
        HIEFFPLA_NET_0_74626);
    
    HIEFFPLA_INST_0_65495 : NOR3B
      port map(A => HIEFFPLA_NET_0_73359, B => 
        HIEFFPLA_NET_0_73276, C => 
        \Science_0/ADC_READ_0/cnt2up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73362);
    
    HIEFFPLA_INST_0_57301 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[43]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75084);
    
    \General_Controller_0/sweep_table_nof_steps[0]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73980, Q => 
        \General_Controller_0/sweep_table_nof_steps[0]_net_1\);
    
    \Timing_0/s_count[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72055, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_count[1]_net_1\);
    
    \Timekeeper_0/microseconds[11]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72149, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[11]\);
    
    HIEFFPLA_INST_0_69868 : AND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72285);
    
    HIEFFPLA_INST_0_69568 : OR3A
      port map(A => HIEFFPLA_NET_0_72410, B => 
        HIEFFPLA_NET_0_72355, C => HIEFFPLA_NET_0_72361, Y => 
        HIEFFPLA_NET_0_72362);
    
    HIEFFPLA_INST_0_62827 : OR3B
      port map(A => HIEFFPLA_NET_0_73969, B => 
        HIEFFPLA_NET_0_73891, C => HIEFFPLA_NET_0_73792, Y => 
        HIEFFPLA_NET_0_73892);
    
    HIEFFPLA_INST_0_59787 : MX2
      port map(A => HIEFFPLA_NET_0_74478, B => 
        HIEFFPLA_NET_0_74570, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74508);
    
    HIEFFPLA_INST_0_57302 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[44]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75083);
    
    \General_Controller_0/sweep_table_samples_per_point[5]\ : 
        DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[5]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[5]_net_1\);
    
    HIEFFPLA_INST_0_68697 : AO1A
      port map(A => HIEFFPLA_NET_0_72668, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_72584);
    
    HIEFFPLA_INST_0_58153 : AO1
      port map(A => \Sensors_0_mag_time[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75145, Y => HIEFFPLA_NET_0_74838);
    
    \General_Controller_0/sweep_table_step_id[5]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73926, Q => 
        \General_Controller_0/sweep_table_step_id[5]_net_1\);
    
    \General_Controller_0/temp_first_byte[3]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73872, Q => 
        \General_Controller_0/temp_first_byte[3]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[12]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[12]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[12]\);
    
    HIEFFPLA_INST_0_70684 : AX1C
      port map(A => \Timing_0/s_time[0]_net_1\, B => 
        HIEFFPLA_NET_0_72058, C => \Timing_0/s_time[1]_net_1\, Y
         => HIEFFPLA_NET_0_72044);
    
    HIEFFPLA_INST_0_64887 : XA1
      port map(A => \I2C_PassThrough_0/cnt[2]_net_1\, B => 
        HIEFFPLA_NET_0_73501, C => HIEFFPLA_NET_0_73515, Y => 
        HIEFFPLA_NET_0_73517);
    
    HIEFFPLA_INST_0_60284 : MX2
      port map(A => \Science_0_chan7_data[0]\, B => 
        \Science_0_chan7_data[4]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74437);
    
    HIEFFPLA_INST_0_65737 : AND2
      port map(A => \Science_0/ADC_READ_0/cnt[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73294);
    
    AFLSDF_INV_36 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_36\);
    
    HIEFFPLA_INST_0_56552 : NOR2A
      port map(A => \Data_Saving_0/Packet_Saver_0/acc_flag_net_1\, 
        B => \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\, Y
         => HIEFFPLA_NET_0_75241);
    
    HIEFFPLA_INST_0_68111 : MX2
      port map(A => HIEFFPLA_NET_0_72726, B => 
        HIEFFPLA_NET_0_72724, S => HIEFFPLA_NET_0_72878, Y => 
        HIEFFPLA_NET_0_72728);
    
    \Science_0/DAC_SET_0/vector[16]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73197, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[16]_net_1\);
    
    HIEFFPLA_INST_0_69871 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_72239, C => HIEFFPLA_NET_0_72227, Y
         => HIEFFPLA_NET_0_72283);
    
    HIEFFPLA_INST_0_60490 : MX2
      port map(A => HIEFFPLA_NET_0_74461, B => 
        HIEFFPLA_NET_0_74477, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74406);
    
    HIEFFPLA_INST_0_62112 : AO1
      port map(A => HIEFFPLA_NET_0_74047, B => 
        HIEFFPLA_NET_0_73900, C => HIEFFPLA_NET_0_74046, Y => 
        HIEFFPLA_NET_0_74050);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_1[10]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74767, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\);
    
    \Science_0/SET_LP_GAIN_0/old_G2[0]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73173, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/old_G2[0]_net_1\);
    
    HIEFFPLA_INST_0_67305 : AO1D
      port map(A => HIEFFPLA_NET_0_72935, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_72736, Y => HIEFFPLA_NET_0_72912);
    
    HIEFFPLA_INST_0_67310 : AO1
      port map(A => HIEFFPLA_NET_0_72935, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        C => HIEFFPLA_NET_0_72924, Y => HIEFFPLA_NET_0_72910);
    
    HIEFFPLA_INST_0_57074 : MX2
      port map(A => HIEFFPLA_NET_0_74944, B => 
        HIEFFPLA_NET_0_74885, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75172);
    
    HIEFFPLA_INST_0_64496 : NOR3B
      port map(A => \General_Controller_0/uc_tx_state[14]_net_1\, 
        B => Communications_0_uc_tx_rdy, C => 
        HIEFFPLA_NET_0_73558, Y => HIEFFPLA_NET_0_73614);
    
    HIEFFPLA_INST_0_71085 : MX2
      port map(A => \GS_Readout_0/state[2]_net_1\, B => 
        \GS_Readout_0/state[1]_net_1\, S => HIEFFPLA_NET_0_74382, 
        Y => HIEFFPLA_NET_0_71981);
    
    HIEFFPLA_INST_0_61687 : MX2
      port map(A => \SweepTable_0_RD[4]\, B => 
        \SweepTable_1_RD[4]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74160);
    
    HIEFFPLA_INST_0_60113 : MX2
      port map(A => \Sensors_0_pressure_raw[18]\, B => 
        \Sensors_0_pressure_raw[22]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74460);
    
    \GS_Readout_0/send[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74714, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74630, Q => 
        \GS_Readout_0_send[3]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[7]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72482, Q => 
        \Sensors_0_gyro_y[7]\);
    
    HIEFFPLA_INST_0_60438 : MX2
      port map(A => \Science_0_chan1_data[11]\, B => 
        \Science_0_chan0_data[3]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74414);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_12\ : DFN1C0
      port map(D => \VCC\, CLK => CLKINT_0_Y_0, CLR => 
        \AFLSDF_INV_7\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_12_Q\);
    
    \Science_0/ADC_READ_0/exp_packet_1[69]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[13]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[69]\);
    
    HIEFFPLA_INST_0_60783 : NOR3B
      port map(A => HIEFFPLA_NET_0_74493, B => 
        HIEFFPLA_NET_0_74433, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74359);
    
    HIEFFPLA_INST_0_57775 : AO1B
      port map(A => \Sensors_0_acc_x[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74945, Y => HIEFFPLA_NET_0_74946);
    
    \Science_0/ADC_READ_0/cnt3dn[6]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73341, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3dn[6]_net_1\);
    
    HIEFFPLA_INST_0_62924 : AOI1D
      port map(A => HIEFFPLA_NET_0_73917, B => 
        HIEFFPLA_NET_0_73904, C => HIEFFPLA_NET_0_73775, Y => 
        HIEFFPLA_NET_0_73865);
    
    HIEFFPLA_INST_0_57239 : AOI1D
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => \Sensors_0_acc_temp[7]\, Y => HIEFFPLA_NET_0_75118);
    
    HIEFFPLA_INST_0_63740 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[2]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[2]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73719);
    
    \ACS_pad/U0/U0\ : IOPAD_TRI
      port map(D => \ACS_pad/U0/NET1\, E => \ACS_pad/U0/NET2\, 
        PAD => ACS);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[11]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72490, Q => 
        \ch3_data_net_0[7]\);
    
    HIEFFPLA_INST_0_61253 : XA1C
      port map(A => 
        \General_Controller_0/state_seconds[13]_net_1\, B => 
        HIEFFPLA_NET_0_74246, C => HIEFFPLA_NET_0_74217, Y => 
        HIEFFPLA_NET_0_74236);
    
    HIEFFPLA_INST_0_70076 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72228);
    
    \Communications_0/FFU_Command_Checker_0/command_out[3]\ : 
        DFN1E1C1
      port map(D => \Communications_0/UART_0_recv[3]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75625, Q => \Communications_0_ext_recv[3]\);
    
    HIEFFPLA_INST_0_57160 : AND2
      port map(A => \Sensors_0_pressure_time[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, Y
         => HIEFFPLA_NET_0_75145);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72335, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\);
    
    \Science_0/ADC_READ_0/g3i[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73257, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73419, Q => 
        \Science_0/ADC_READ_0_G3[0]\);
    
    HIEFFPLA_INST_0_69043 : NAND2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        B => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72488);
    
    HIEFFPLA_INST_0_69134 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[6]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[7]_net_1\, 
        C => HIEFFPLA_NET_0_72556, Y => HIEFFPLA_NET_0_72463);
    
    HIEFFPLA_INST_0_71132 : AOI1D
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => \Sensors_0_acc_temp[3]\, Y => HIEFFPLA_NET_0_71976);
    
    HIEFFPLA_INST_0_62203 : AND3B
      port map(A => CLKINT_1_Y, B => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, C => 
        HIEFFPLA_NET_0_74030, Y => HIEFFPLA_NET_0_74031);
    
    HIEFFPLA_INST_0_55046 : AND2
      port map(A => HIEFFPLA_NET_0_75593, B => 
        HIEFFPLA_NET_0_75591, Y => HIEFFPLA_NET_0_75604);
    
    \Science_0/ADC_READ_0/cnt1dn[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73408, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1dn[0]_net_1\);
    
    \General_Controller_0/sweep_table_samples_per_point[7]\ : 
        DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[7]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[7]_net_1\);
    
    HIEFFPLA_INST_0_55723 : AO1
      port map(A => HIEFFPLA_NET_0_75438, B => 
        \Communications_0/UART_1/rx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_75433, Y => HIEFFPLA_NET_0_75437);
    
    \Data_Saving_0/Packet_Saver_0/old_acc_new_data\ : DFN0P1
      port map(D => \AFLSDF_INV_8\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => 
        \Data_Saving_0/Packet_Saver_0/old_acc_new_data_i_0\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/data_out[2]\ : DFN0E1C1
      port map(D => GYRO_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72681, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[2]\);
    
    \Science_0/DAC_SET_0/vector[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73194, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[2]_net_1\);
    
    HIEFFPLA_INST_0_68583 : AO1A
      port map(A => HIEFFPLA_NET_0_72602, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\, C
         => \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_72612);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[0]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72754, Q => 
        \Sensors_0_acc_z[0]\);
    
    HIEFFPLA_INST_0_69063 : NOR3B
      port map(A => HIEFFPLA_NET_0_72492, B => 
        HIEFFPLA_NET_0_72540, C => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_72480);
    
    HIEFFPLA_INST_0_57139 : AND2
      port map(A => \Sensors_0_pressure_temp_raw[19]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75158);
    
    \General_Controller_0/uc_pwr_en\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74120, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => UC_PWR_EN_c);
    
    HIEFFPLA_INST_0_62831 : XNOR2
      port map(A => \General_Controller_0/uc_rx_state[3]_net_1\, 
        B => \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73890);
    
    HIEFFPLA_INST_0_70880 : NAND3C
      port map(A => HIEFFPLA_NET_0_72006, B => 
        HIEFFPLA_NET_0_72796, C => HIEFFPLA_NET_0_72781, Y => 
        HIEFFPLA_NET_0_72748);
    
    \Science_0/ADC_READ_0/data_a[7]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[7]_net_1\);
    
    HIEFFPLA_INST_0_58214 : AND2
      port map(A => \Sensors_0_acc_y[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        Y => HIEFFPLA_NET_0_74826);
    
    HIEFFPLA_INST_0_61984 : XA1
      port map(A => \General_Controller_0/uc_rx_byte[4]_net_1\, B
         => \General_Controller_0/uc_rx_byte[2]_net_1\, C => 
        HIEFFPLA_NET_0_73803, Y => HIEFFPLA_NET_0_74083);
    
    \L1WR_pad/U0/U0\ : IOPAD_TRI
      port map(D => \L1WR_pad/U0/NET1\, E => \L1WR_pad/U0/NET2\, 
        PAD => L1WR);
    
    HIEFFPLA_INST_0_59497 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[1]\, B => 
        \Data_Hub_Packets_0_status_packet[5]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74546);
    
    HIEFFPLA_INST_0_65660 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt4dn[3]_net_1\, B => 
        HIEFFPLA_NET_0_73329, C => HIEFFPLA_NET_0_73274, Y => 
        HIEFFPLA_NET_0_73315);
    
    \General_Controller_0/sweep_table_probe_id[3]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73924, Q => 
        \General_Controller_0/sweep_table_probe_id[3]_net_1\);
    
    \Science_0/ADC_READ_0/data_a[1]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[0]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[1]_net_1\);
    
    HIEFFPLA_INST_0_69587 : AOI1D
      port map(A => HIEFFPLA_NET_0_72426, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72358);
    
    HIEFFPLA_INST_0_59955 : MX2
      port map(A => \Sensors_0_pressure_raw[16]\, B => 
        \Sensors_0_pressure_raw[20]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74483);
    
    HIEFFPLA_INST_0_57687 : AO1B
      port map(A => \Sensors_0_gyro_y[13]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74969, Y => HIEFFPLA_NET_0_74970);
    
    HIEFFPLA_INST_0_55980 : NAND2B
      port map(A => UC_UART_TX_c, B => UC_CONSOLE_EN_c, Y => 
        HIEFFPLA_NET_0_75378);
    
    \Data_Saving_0/Packet_Saver_0/data_out[7]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75206, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[7]\);
    
    \Pressure_Signal_Debounce_0/ms_cnt[1]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73494, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[1]_net_1\);
    
    HIEFFPLA_INST_0_68501 : OR2A
      port map(A => HIEFFPLA_NET_0_72619, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_net_1\, Y => 
        HIEFFPLA_NET_0_72635);
    
    HIEFFPLA_INST_0_57557 : AND2
      port map(A => \Sensors_0_gyro_time[19]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75010);
    
    \Science_0/DAC_SET_0/sdi_int\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73214, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73213, Q => 
        LDSDI_c);
    
    HIEFFPLA_INST_0_61936 : NOR3B
      port map(A => \General_Controller_0/uc_rx_byte[7]_net_1\, B
         => \General_Controller_0/uc_rx_substate[2]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74094);
    
    HIEFFPLA_INST_0_59621 : MX2
      port map(A => \Sensors_0_pressure_temp_raw[21]\, B => 
        \Sensors_0_pressure_raw[13]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74530);
    
    HIEFFPLA_INST_0_70149 : AO1C
      port map(A => \Sensors_0/Pressure_Sensor_0/state[8]\, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]_net_1\, 
        C => HIEFFPLA_NET_0_72241, Y => HIEFFPLA_NET_0_72209);
    
    HIEFFPLA_INST_0_60431 : NOR3B
      port map(A => HIEFFPLA_NET_0_74415, B => 
        HIEFFPLA_NET_0_74341, C => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74416);
    
    HIEFFPLA_INST_0_59557 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[48]\, B => 
        \Data_Hub_Packets_0_status_packet[52]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74538);
    
    HIEFFPLA_INST_0_67140 : NOR3A
      port map(A => HIEFFPLA_NET_0_72955, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[3]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72954);
    
    HIEFFPLA_INST_0_63042 : AOI1
      port map(A => \General_Controller_0/uc_rx_byte[4]_net_1\, B
         => \General_Controller_0/uc_rx_byte[0]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73842);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[3]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72808, Q => 
        \Sensors_0_mag_z[3]\);
    
    HIEFFPLA_INST_0_60528 : AO1
      port map(A => HIEFFPLA_NET_0_74541, B => 
        HIEFFPLA_NET_0_74341, C => HIEFFPLA_NET_0_74400, Y => 
        HIEFFPLA_NET_0_74401);
    
    HIEFFPLA_INST_0_57392 : AO1
      port map(A => \Sensors_0_gyro_temp[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75057, Y => HIEFFPLA_NET_0_75058);
    
    \General_Controller_0/constant_bias_probe_id[2]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73923, Q => 
        \General_Controller_0/un10_uc_tx_rdy_i[2]\);
    
    \FRAM_SDA_pad/U0/U1\ : IOBI_IB_OB_EB
      port map(D => \GND\, E => \I2C_PassThrough_0.state[3]\, YIN
         => \FRAM_SDA_pad/U0/NET3\, DOUT => 
        \FRAM_SDA_pad/U0/NET1\, EOUT => \FRAM_SDA_pad/U0/NET2\, Y
         => FRAM_SDA_in);
    
    HIEFFPLA_INST_0_57621 : AO1
      port map(A => \Sensors_0_pressure_raw[15]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74989, Y => HIEFFPLA_NET_0_74990);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[5]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[5]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[5]\);
    
    HIEFFPLA_INST_0_63140 : AO1
      port map(A => HIEFFPLA_NET_0_73930, B => 
        \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        HIEFFPLA_NET_0_73843, Y => HIEFFPLA_NET_0_73821);
    
    HIEFFPLA_INST_0_66447 : AND3
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        B => ACCE_SCL_c, C => HIEFFPLA_NET_0_73118, Y => 
        HIEFFPLA_NET_0_73119);
    
    HIEFFPLA_INST_0_67372 : AO1
      port map(A => HIEFFPLA_NET_0_72918, B => 
        HIEFFPLA_NET_0_72760, C => HIEFFPLA_NET_0_72887, Y => 
        HIEFFPLA_NET_0_72896);
    
    HIEFFPLA_INST_0_57697 : AO1B
      port map(A => \Sensors_0_acc_y[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74966, Y => HIEFFPLA_NET_0_74967);
    
    HIEFFPLA_INST_0_68954 : NOR2A
      port map(A => HIEFFPLA_NET_0_72543, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, Y
         => HIEFFPLA_NET_0_72514);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[5]\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72295, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72221, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[5]_net_1\);
    
    HIEFFPLA_INST_0_65951 : NAND3A
      port map(A => HIEFFPLA_NET_0_73350, B => 
        \Science_0/ADC_READ_0/cnt3up[4]_net_1\, C => 
        HIEFFPLA_NET_0_73276, Y => HIEFFPLA_NET_0_73253);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[1]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[1]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[1]\);
    
    HIEFFPLA_INST_0_66179 : MX2B
      port map(A => \Science_0/DAC_SET_0/vector[8]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73187);
    
    HIEFFPLA_INST_0_61620 : NOR2A
      port map(A => HIEFFPLA_NET_0_74181, B => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74172);
    
    HIEFFPLA_INST_0_67551 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        B => HIEFFPLA_NET_0_72741, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, Y
         => HIEFFPLA_NET_0_72854);
    
    HIEFFPLA_INST_0_62037 : NAND3C
      port map(A => HIEFFPLA_NET_0_74064, B => 
        HIEFFPLA_NET_0_74061, C => HIEFFPLA_NET_0_74090, Y => 
        HIEFFPLA_NET_0_74065);
    
    HIEFFPLA_INST_0_55117 : AO1C
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[28]_net_1\, B => 
        HIEFFPLA_NET_0_75578, C => 
        \Communications_0/UART_0/rx_clk_count[27]_net_1\, Y => 
        HIEFFPLA_NET_0_75585);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[18]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[18]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[18]\);
    
    HIEFFPLA_INST_0_57837 : AO1B
      port map(A => \Sensors_0_mag_time[19]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74929, Y => HIEFFPLA_NET_0_74930);
    
    \General_Controller_0/sweep_table_sweep_cnt[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74144, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[0]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRYSYNC[7]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_7_Q\, CLK
         => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[7]\\\\\);
    
    \Science_0/ADC_READ_0/cnt3dn[4]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73343, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3dn[4]_net_1\);
    
    HIEFFPLA_INST_0_71131 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_71976, Y => HIEFFPLA_NET_0_75073);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[4]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_75249, CLK => CLKINT_0_Y_0, E
         => CLKINT_1_Y, Q => 
        \Data_Saving_0/Interrupt_Generator_0/counter[4]_net_1\);
    
    \Science_0/ADC_READ_0/chan2_data[1]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[1]\);
    
    HIEFFPLA_INST_0_62318 : OA1C
      port map(A => Communications_0_uc_rx_rdy, B => 
        \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        HIEFFPLA_NET_0_74006, Y => HIEFFPLA_NET_0_74007);
    
    \GS_Readout_0/subState_RNITID3[0]\ : CLKINT
      port map(A => \GS_Readout_0/subState_0[0]\, Y => 
        \GS_Readout_0/subState[0]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[6]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72783, Q => 
        \Sensors_0_mag_y[6]\);
    
    HIEFFPLA_INST_0_55977 : MX2
      port map(A => \Communications_0/UART_0_tx\, B => 
        UC_UART_TX_c, S => UC_CONSOLE_EN_c, Y => SCIENCE_TX_c_c);
    
    \General_Controller_0/sweep_table_points[9]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[9]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72266, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\);
    
    \General_Controller_0/uc_tx_state[7]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73566, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[7]_net_1\);
    
    \FMC_DA_pad[1]/U0/U0\ : IOPAD_TRI
      port map(D => \FMC_DA_pad[1]/U0/NET1\, E => 
        \FMC_DA_pad[1]/U0/NET2\, PAD => FMC_DA(1));
    
    HIEFFPLA_INST_0_63526 : MX2
      port map(A => HIEFFPLA_NET_0_73679, B => 
        HIEFFPLA_NET_0_73671, S => HIEFFPLA_NET_0_73621, Y => 
        HIEFFPLA_NET_0_73754);
    
    HIEFFPLA_INST_0_57314 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_75078, Y => HIEFFPLA_NET_0_75079);
    
    HIEFFPLA_INST_0_56424 : MX2
      port map(A => \FMC_DA_c[3]\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[3]\\\\\, S => 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\, Y => 
        HIEFFPLA_NET_0_75284);
    
    \Science_0/ADC_READ_0/g1i[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73266, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0_G1[0]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[21]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72282, Q => 
        \Sensors_0_pressure_temp_raw[21]\);
    
    \Science_0/ADC_READ_0/cnt1dn[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73406, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1dn[2]_net_1\);
    
    HIEFFPLA_INST_0_68520 : NOR2A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[2]_net_1\, B => 
        HIEFFPLA_NET_0_72705, Y => HIEFFPLA_NET_0_72629);
    
    \General_Controller_0/uc_tx_nextstate[4]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73973, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73857, Q => 
        \General_Controller_0/uc_tx_nextstate[4]_net_1\);
    
    HIEFFPLA_INST_0_69697 : AOI1D
      port map(A => HIEFFPLA_NET_0_72346, B => 
        HIEFFPLA_NET_0_72424, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72326);
    
    HIEFFPLA_INST_0_56662 : MX2
      port map(A => HIEFFPLA_NET_0_75194, B => 
        HIEFFPLA_NET_0_75058, S => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75227);
    
    HIEFFPLA_INST_0_64749 : MX2
      port map(A => HIEFFPLA_NET_0_73614, B => 
        HIEFFPLA_NET_0_73530, S => HIEFFPLA_NET_0_73521, Y => 
        HIEFFPLA_NET_0_73549);
    
    HIEFFPLA_INST_0_69922 : AO1
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[1]_net_1\, 
        B => HIEFFPLA_NET_0_72238, C => HIEFFPLA_NET_0_72260, Y
         => HIEFFPLA_NET_0_72266);
    
    HIEFFPLA_INST_0_60996 : AND2
      port map(A => \General_Controller_0/ext_rx_state_i_0[1]\, B
         => Communications_0_ext_rx_rdy, Y => 
        HIEFFPLA_NET_0_74301);
    
    HIEFFPLA_INST_0_67826 : AND3
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => \Sensors_0/Accelerometer_0/state_0[8]\, Y => 
        HIEFFPLA_NET_0_72793);
    
    \General_Controller_0/uc_tx_substate[3]\ : DFN1C1
      port map(D => 
        \General_Controller_0/uc_tx_substate[3]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_tx_substate[3]_net_1\);
    
    HIEFFPLA_INST_0_60023 : MX2
      port map(A => HIEFFPLA_NET_0_74566, B => 
        HIEFFPLA_NET_0_74446, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74472);
    
    HIEFFPLA_INST_0_57742 : NAND3C
      port map(A => HIEFFPLA_NET_0_74840, B => 
        HIEFFPLA_NET_0_74832, C => HIEFFPLA_NET_0_74817, Y => 
        HIEFFPLA_NET_0_74955);
    
    HIEFFPLA_INST_0_57272 : AND2
      port map(A => \ch3_data_net_0[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75099);
    
    HIEFFPLA_INST_0_69897 : AND2B
      port map(A => HIEFFPLA_NET_0_72278, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72274);
    
    HIEFFPLA_INST_0_58552 : XNOR2
      port map(A => FFU_EJECTED_c, B => 
        \Eject_Signal_Debounce_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74736);
    
    HIEFFPLA_INST_0_57412 : AO1
      port map(A => \ch3_data_net_0[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74875, Y => HIEFFPLA_NET_0_75053);
    
    HIEFFPLA_INST_0_70626 : NAND3B
      port map(A => \Timing_0/s_count[2]_net_1\, B => 
        \Timing_0/s_count[0]_net_1\, C => 
        \Timing_0/s_count[6]_net_1\, Y => HIEFFPLA_NET_0_72060);
    
    HIEFFPLA_INST_0_59033 : NOR3B
      port map(A => HIEFFPLA_NET_0_74507, B => 
        HIEFFPLA_NET_0_74649, C => HIEFFPLA_NET_0_74574, Y => 
        HIEFFPLA_NET_0_74631);
    
    HIEFFPLA_INST_0_63128 : AO1A
      port map(A => HIEFFPLA_NET_0_73847, B => 
        HIEFFPLA_NET_0_74094, C => HIEFFPLA_NET_0_73846, Y => 
        HIEFFPLA_NET_0_73823);
    
    HIEFFPLA_INST_0_58158 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[12]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75144, Y => HIEFFPLA_NET_0_74837);
    
    HIEFFPLA_INST_0_57054 : AOI1D
      port map(A => HIEFFPLA_NET_0_74838, B => 
        HIEFFPLA_NET_0_74949, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75175);
    
    HIEFFPLA_INST_0_56538 : AX1C
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[5]_net_1\, B
         => HIEFFPLA_NET_0_75254, C => 
        \Data_Saving_0/Interrupt_Generator_0/counter[6]_net_1\, Y
         => HIEFFPLA_NET_0_75247);
    
    HIEFFPLA_INST_0_61905 : AND3
      port map(A => HIEFFPLA_NET_0_73803, B => 
        HIEFFPLA_NET_0_74101, C => HIEFFPLA_NET_0_74091, Y => 
        HIEFFPLA_NET_0_74102);
    
    HIEFFPLA_INST_0_63560 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[12]_net_1\, B
         => \General_Controller_0/sweep_table_points[12]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73749);
    
    HIEFFPLA_INST_0_68783 : NAND2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        B => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72563);
    
    \LDCS_pad/U0/U0\ : IOPAD_TRI
      port map(D => \LDCS_pad/U0/NET1\, E => \LDCS_pad/U0/NET2\, 
        PAD => LDCS);
    
    HIEFFPLA_INST_0_60213 : MX2
      port map(A => HIEFFPLA_NET_0_74479, B => 
        HIEFFPLA_NET_0_74503, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74445);
    
    \Communications_0/FFU_Command_Checker_0/command_out[6]\ : 
        DFN1E1C1
      port map(D => \Communications_0/UART_0_recv[6]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75625, Q => \Communications_0_ext_recv[6]\);
    
    HIEFFPLA_INST_0_56114 : XO1A
      port map(A => HIEFFPLA_NET_0_75366, B => 
        HIEFFPLA_NET_0_89701, C => HIEFFPLA_NET_0_75343, Y => 
        HIEFFPLA_NET_0_75344);
    
    \Science_0/ADC_READ_0/chan3_data[10]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[10]\);
    
    HIEFFPLA_INST_0_70971 : OR3B
      port map(A => HIEFFPLA_NET_0_73054, B => 
        HIEFFPLA_NET_0_73010, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_71998);
    
    \I2C_PassThrough_0/cnt[3]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73502, CLK => CLKINT_0_Y_0, Q
         => \I2C_PassThrough_0/cnt[3]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[19]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72282, Q => 
        \Sensors_0_pressure_temp_raw[19]\);
    
    \Science_0/ADC_READ_0/data_a[13]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[13]_net_1\);
    
    HIEFFPLA_INST_0_60373 : MX2
      port map(A => \Science_0_chan1_data[10]\, B => 
        \Science_0_chan0_data[2]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74425);
    
    \General_Controller_0/sweep_table_sweep_cnt[13]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74140, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[13]_net_1\);
    
    HIEFFPLA_INST_0_70548 : AND2
      port map(A => HIEFFPLA_NET_0_72082, B => 
        HIEFFPLA_NET_0_72081, Y => HIEFFPLA_NET_0_72083);
    
    \Communications_0/UART_0/rx_clk_count[24]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75575, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75554, Q => 
        \Communications_0/UART_0/rx_clk_count[24]_net_1\);
    
    HIEFFPLA_INST_0_66584 : MX2
      port map(A => HIEFFPLA_NET_0_73085, B => 
        HIEFFPLA_NET_0_73084, S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73088);
    
    HIEFFPLA_INST_0_66303 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[0]\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73150);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_13\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[7]\\\\\, CLK => 
        CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_13_Q\);
    
    HIEFFPLA_INST_0_56564 : MX2
      port map(A => HIEFFPLA_NET_0_75237, B => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, S => 
        \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\, Y => 
        HIEFFPLA_NET_0_75238);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[1]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72801, Q => 
        \Sensors_0_acc_x[1]\);
    
    HIEFFPLA_INST_0_69588 : AND2
      port map(A => HIEFFPLA_NET_0_72410, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72357);
    
    HIEFFPLA_INST_0_61996 : AND3
      port map(A => HIEFFPLA_NET_0_74087, B => 
        \General_Controller_0/uc_rx_byte[1]_net_1\, C => 
        HIEFFPLA_NET_0_73881, Y => HIEFFPLA_NET_0_74078);
    
    HIEFFPLA_INST_0_56328 : XOR2
      port map(A => HIEFFPLA_NET_0_75291, B => 
        HIEFFPLA_NET_0_75288, Y => HIEFFPLA_NET_0_75309);
    
    HIEFFPLA_INST_0_69444 : AND2
      port map(A => HIEFFPLA_NET_0_72430, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_i2c_addr[0]\, 
        Y => HIEFFPLA_NET_0_72387);
    
    HIEFFPLA_INST_0_69306 : OR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72423);
    
    HIEFFPLA_INST_0_66265 : MX2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G4[1]_net_1\, B
         => \Science_0/ADC_READ_0_G4[1]\, S => 
        \Science_0/SET_LP_GAIN_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73162);
    
    HIEFFPLA_INST_0_65400 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt1up[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt1up[0]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt1up[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73388);
    
    HIEFFPLA_INST_0_70188 : NAND3B
      port map(A => HIEFFPLA_NET_0_72311, B => 
        HIEFFPLA_NET_0_72198, C => 
        \Sensors_0/Pressure_Sensor_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72199);
    
    HIEFFPLA_INST_0_59300 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[50]\, B => 
        \Data_Hub_Packets_0_status_packet[54]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74572);
    
    HIEFFPLA_INST_0_57730 : NAND3C
      port map(A => HIEFFPLA_NET_0_74842, B => 
        HIEFFPLA_NET_0_74833, C => HIEFFPLA_NET_0_74819, Y => 
        HIEFFPLA_NET_0_74958);
    
    HIEFFPLA_INST_0_66017 : AND3C
      port map(A => \Science_0/ADC_READ_0/state[2]_net_1\, B => 
        \Science_0/ADC_READ_0/state[1]_net_1\, C => 
        HIEFFPLA_NET_0_73239, Y => HIEFFPLA_NET_0_73237);
    
    HIEFFPLA_INST_0_64101 : MX2
      port map(A => HIEFFPLA_NET_0_73634, B => 
        HIEFFPLA_NET_0_73626, S => HIEFFPLA_NET_0_73585, Y => 
        HIEFFPLA_NET_0_73671);
    
    HIEFFPLA_INST_0_55075 : AND3C
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[29]_net_1\, B => 
        \Communications_0/UART_0/rx_clk_count[30]_net_1\, C => 
        \Communications_0/UART_0/rx_clk_count_c0\, Y => 
        HIEFFPLA_NET_0_75597);
    
    HIEFFPLA_INST_0_64850 : AO1C
      port map(A => HIEFFPLA_NET_0_73560, B => 
        HIEFFPLA_NET_0_73597, C => HIEFFPLA_NET_0_73524, Y => 
        HIEFFPLA_NET_0_73525);
    
    HIEFFPLA_INST_0_57333 : AOI1
      port map(A => \Science_0_exp_packet_0[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_75073, Y => HIEFFPLA_NET_0_75074);
    
    \General_Controller_0/st_wdata[12]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[12]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[12]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[8]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72807, Q => 
        \Sensors_0_mag_z[8]\);
    
    HIEFFPLA_INST_0_61870 : OR3B
      port map(A => HIEFFPLA_NET_0_74094, B => 
        \General_Controller_0/uc_rx_byte[3]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74112);
    
    \General_Controller_0/sweep_table_samples_per_step[3]\ : 
        DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[3]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[3]_net_1\);
    
    \Timekeeper_0/milliseconds[10]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72115, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[10]\);
    
    \General_Controller_0/sweep_table_samples_per_step[14]\ : 
        DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[14]_net_1\);
    
    HIEFFPLA_INST_0_67351 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        C => HIEFFPLA_NET_0_72929, Y => HIEFFPLA_NET_0_72901);
    
    HIEFFPLA_INST_0_62385 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state_0[3]_net_1\, 
        B => \General_Controller_0/uc_rx_substate[2]_net_1\, C
         => \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73992);
    
    HIEFFPLA_INST_0_71065 : AO1A
      port map(A => \GS_Readout_0/prevState[0]_net_1\, B => 
        HIEFFPLA_NET_0_71983, C => HIEFFPLA_NET_0_74587, Y => 
        HIEFFPLA_NET_0_74598);
    
    \Communications_0/UART_1/tx_clk_count[6]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75405, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_clk_count_i_0[6]\);
    
    \Science_0/DAC_SET_0/vector[15]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73198, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[15]_net_1\);
    
    HIEFFPLA_INST_0_66546 : OR3A
      port map(A => HIEFFPLA_NET_0_73045, B => 
        HIEFFPLA_NET_0_73093, C => HIEFFPLA_NET_0_73092, Y => 
        HIEFFPLA_NET_0_73094);
    
    \General_Controller_0/uc_rx_byte_0[2]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[2]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte_0[2]_net_1\);
    
    \General_Controller_0/status_bits_1[43]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74203, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[43]\);
    
    HIEFFPLA_INST_0_69351 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[2]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72411);
    
    HIEFFPLA_INST_0_64217 : MX2
      port map(A => HIEFFPLA_NET_0_73744, B => 
        HIEFFPLA_NET_0_73736, S => HIEFFPLA_NET_0_73588, Y => 
        HIEFFPLA_NET_0_73648);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[3]\ : 
        DFN1E1
      port map(D => CLKINT_1_Y, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_72919, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[3]_net_1\);
    
    HIEFFPLA_INST_0_70543 : AX1C
      port map(A => HIEFFPLA_NET_0_72090, B => 
        \Timing_0/f_time[3]_net_1\, C => \s_clks_net_0[4]\, Y => 
        HIEFFPLA_NET_0_72086);
    
    HIEFFPLA_INST_0_67734 : AND3A
      port map(A => HIEFFPLA_NET_0_72914, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        C => \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        Y => HIEFFPLA_NET_0_72813);
    
    HIEFFPLA_INST_0_66187 : AOI1
      port map(A => \Science_0/SET_LP_GAIN_0/state[7]_net_1\, B
         => \Science_0/ADC_READ_0_G1[0]\, C => 
        HIEFFPLA_NET_0_73183, Y => HIEFFPLA_NET_0_73184);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[2]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72276, Q => \Sensors_0_pressure_raw[2]\);
    
    HIEFFPLA_INST_0_65320 : NOR3B
      port map(A => \Science_0/ADC_READ_0/cnt1dn[3]_net_1\, B => 
        HIEFFPLA_NET_0_73411, C => 
        \Science_0/ADC_READ_0/cnt1dn[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73412);
    
    HIEFFPLA_INST_0_56370 : AX1A
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, B
         => HIEFFPLA_NET_0_75370, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, Y
         => HIEFFPLA_NET_0_75298);
    
    HIEFFPLA_INST_0_55456 : AO1
      port map(A => HIEFFPLA_NET_0_75512, B => 
        \Communications_0/UART_0/tx_count[1]_net_1\, C => 
        HIEFFPLA_NET_0_75506, Y => HIEFFPLA_NET_0_75507);
    
    HIEFFPLA_INST_0_58626 : AO1D
      port map(A => HIEFFPLA_NET_0_74707, B => 
        HIEFFPLA_NET_0_74655, C => HIEFFPLA_NET_0_74691, Y => 
        HIEFFPLA_NET_0_74717);
    
    HIEFFPLA_INST_0_69021 : NOR2A
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72495);
    
    HIEFFPLA_INST_0_61295 : AX1B
      port map(A => HIEFFPLA_NET_0_74217, B => 
        HIEFFPLA_NET_0_74262, C => HIEFFPLA_NET_0_74224, Y => 
        HIEFFPLA_NET_0_74225);
    
    \Science_0/DAC_SET_0/vector[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73191, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[5]_net_1\);
    
    HIEFFPLA_INST_0_70396 : AX1C
      port map(A => \Timekeeper_0_microseconds[9]\, B => 
        HIEFFPLA_NET_0_72157, C => 
        \Timekeeper_0_microseconds[10]\, Y => 
        HIEFFPLA_NET_0_72150);
    
    \GYRO_SDA_pad/U0/U0\ : IOPAD_BI
      port map(D => \GYRO_SDA_pad/U0/NET1\, E => 
        \GYRO_SDA_pad/U0/NET2\, Y => \GYRO_SDA_pad/U0/NET3\, PAD
         => GYRO_SDA);
    
    HIEFFPLA_INST_0_58066 : AO1
      port map(A => \Sensors_0_gyro_y[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75158, Y => HIEFFPLA_NET_0_74865);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72262, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\);
    
    \Timekeeper_0/milliseconds[8]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72094, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[8]\);
    
    HIEFFPLA_INST_0_60862 : NAND2B
      port map(A => HIEFFPLA_NET_0_74328, B => 
        HIEFFPLA_NET_0_74330, Y => HIEFFPLA_NET_0_74337);
    
    HIEFFPLA_INST_0_55243 : AND2B
      port map(A => \Communications_0/UART_0/rx_state[0]_net_1\, 
        B => \Communications_0/UART_0/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75554);
    
    HIEFFPLA_INST_0_70091 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72222);
    
    HIEFFPLA_INST_0_64702 : OR3A
      port map(A => 
        \General_Controller_0/uc_tx_substate[2]_net_1\, B => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, C => 
        HIEFFPLA_NET_0_73563, Y => HIEFFPLA_NET_0_73559);
    
    HIEFFPLA_INST_0_59885 : MX2
      port map(A => \Science_0_chan1_data[2]\, B => 
        \Science_0_chan1_data[6]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74492);
    
    HIEFFPLA_INST_0_62211 : AND2
      port map(A => HIEFFPLA_NET_0_74027, B => 
        HIEFFPLA_NET_0_73778, Y => HIEFFPLA_NET_0_74028);
    
    \Data_Saving_0/Packet_Saver_0/packet_select[11]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74772, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\);
    
    HIEFFPLA_INST_0_68760 : NAND3C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, C
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72568);
    
    HIEFFPLA_INST_0_54934 : NOR3B
      port map(A => \ClockDivs_0/cnt_800kHz[4]_net_1\, B => 
        \ClockDivs_0/cnt_800kHz[0]_net_1\, C => 
        \ClockDivs_0/cnt_800kHz[3]_net_1\, Y => 
        HIEFFPLA_NET_0_75635);
    
    AFLSDF_INV_9 : INV
      port map(A => \Timing_0/f_time[0]_net_1\, Y => 
        \AFLSDF_INV_9\);
    
    HIEFFPLA_INST_0_57387 : AO1
      port map(A => \Data_Hub_Packets_0_status_packet[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, C
         => HIEFFPLA_NET_0_75059, Y => HIEFFPLA_NET_0_75060);
    
    \General_Controller_0/sweep_table_write_value[2]\ : DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[2]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[2]_net_1\);
    
    \Communications_0/UART_0/recv[0]\ : DFN1E1C1
      port map(D => \Communications_0/UART_0/rx_byte[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75551, Q => 
        \Communications_0/UART_0_recv[0]\);
    
    HIEFFPLA_INST_0_62667 : AND3
      port map(A => HIEFFPLA_NET_0_73958, B => 
        HIEFFPLA_NET_0_73775, C => 
        \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73932);
    
    HIEFFPLA_INST_0_58439 : NOR3A
      port map(A => HIEFFPLA_NET_0_74771, B => 
        \Data_Saving_0/Packet_Saver_0/gyro_flag_net_1\, C => 
        \Data_Saving_0/Packet_Saver_0/pressure_flag_net_1\, Y => 
        HIEFFPLA_NET_0_74766);
    
    HIEFFPLA_INST_0_69938 : AO1D
      port map(A => HIEFFPLA_NET_0_72257, B => 
        HIEFFPLA_NET_0_72238, C => HIEFFPLA_NET_0_72252, Y => 
        HIEFFPLA_NET_0_72263);
    
    \Science_0/ADC_READ_0/cnt3up[3]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73333, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3up[3]_net_1\);
    
    HIEFFPLA_INST_0_61622 : NOR2A
      port map(A => HIEFFPLA_NET_0_74181, B => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_74171);
    
    HIEFFPLA_INST_0_59509 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[43]\, B => 
        \Data_Hub_Packets_0_status_packet[47]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74544);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[2]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[2]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[2]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[4]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72489, Q => 
        \ch3_data_net_0[0]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[5]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72804, Q => 
        \Sensors_0_mag_x[5]\);
    
    HIEFFPLA_INST_0_66626 : AND3A
      port map(A => ACCE_SCL_c, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        C => HIEFFPLA_NET_0_73090, Y => HIEFFPLA_NET_0_73079);
    
    HIEFFPLA_INST_0_64715 : AOI1C
      port map(A => \General_Controller_0/uc_tx_state[5]_net_1\, 
        B => \General_Controller_0/uc_tx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_73559, Y => HIEFFPLA_NET_0_73554);
    
    HIEFFPLA_INST_0_64677 : AND2
      port map(A => 
        \General_Controller_0/uc_tx_nextstate[6]_net_1\, B => 
        HIEFFPLA_NET_0_73584, Y => HIEFFPLA_NET_0_73567);
    
    \General_Controller_0/uc_rx_substate[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73771, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_substate[3]_net_1\);
    
    HIEFFPLA_INST_0_64675 : AND2
      port map(A => 
        \General_Controller_0/uc_tx_nextstate[5]_net_1\, B => 
        HIEFFPLA_NET_0_73584, Y => HIEFFPLA_NET_0_73568);
    
    HIEFFPLA_INST_0_63999 : MX2
      port map(A => HIEFFPLA_NET_0_73652, B => 
        HIEFFPLA_NET_0_73644, S => HIEFFPLA_NET_0_73599, Y => 
        HIEFFPLA_NET_0_73681);
    
    HIEFFPLA_INST_0_69647 : OA1C
      port map(A => HIEFFPLA_NET_0_72330, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[2]_net_1\, 
        C => HIEFFPLA_NET_0_72325, Y => HIEFFPLA_NET_0_72337);
    
    HIEFFPLA_INST_0_66953 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        B => \Sensors_0/Accelerometer_0/state_0[8]\, C => 
        HIEFFPLA_NET_0_72799, Y => HIEFFPLA_NET_0_72997);
    
    HIEFFPLA_INST_0_58783 : NAND3C
      port map(A => HIEFFPLA_NET_0_74700, B => 
        HIEFFPLA_NET_0_74673, C => HIEFFPLA_NET_0_74685, Y => 
        HIEFFPLA_NET_0_74686);
    
    HIEFFPLA_INST_0_66563 : AO1
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        B => ACCE_SCL_c, C => HIEFFPLA_NET_0_73047, Y => 
        HIEFFPLA_NET_0_73091);
    
    \Communications_0/FFU_Command_Checker_0/state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75622, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/FFU_Command_Checker_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_57920 : AOI1
      port map(A => \Sensors_0_acc_time[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74904, Y => HIEFFPLA_NET_0_74905);
    
    \Communications_0/UART_0/recv[2]\ : DFN1E1C1
      port map(D => \Communications_0/UART_0/rx_byte[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75551, Q => 
        \Communications_0/UART_0_recv[2]\);
    
    HIEFFPLA_INST_0_65519 : NAND2B
      port map(A => \Science_0/ADC_READ_0/cnt3dn[2]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt3dn[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73355);
    
    HIEFFPLA_INST_0_62498 : NOR2A
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => CLKINT_1_Y, Y => HIEFFPLA_NET_0_73970);
    
    HIEFFPLA_INST_0_55276 : MX2A
      port map(A => HIEFFPLA_NET_0_75380, B => 
        HIEFFPLA_NET_0_75583, S => 
        \Communications_0/UART_0/rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75547);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/sda_1\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_73094, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73064, Q => 
        \Sensors_0.Accelerometer_0.I2C_Master_0.sda_1\);
    
    HIEFFPLA_INST_0_64129 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_1[9]_net_1\, 
        B => 
        \General_Controller_0/constant_bias_voltage_1[1]_net_1\, 
        S => HIEFFPLA_NET_0_73558, Y => HIEFFPLA_NET_0_73664);
    
    \General_Controller_0/uc_rx_byte[4]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[4]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte[4]_net_1\);
    
    \Pressure_Signal_Debounce_0/ms_cnt[9]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73484, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[9]_net_1\);
    
    \General_Controller_0/constant_bias_voltage_1[10]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[10]_net_1\);
    
    HIEFFPLA_INST_0_68980 : NOR3A
      port map(A => HIEFFPLA_NET_0_72507, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[7]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72508);
    
    HIEFFPLA_INST_0_66761 : NAND3C
      port map(A => HIEFFPLA_NET_0_73050, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        C => HIEFFPLA_NET_0_73051, Y => HIEFFPLA_NET_0_73041);
    
    HIEFFPLA_INST_0_66134 : MX2B
      port map(A => \Science_0/DAC_SET_0/vector[14]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73198);
    
    HIEFFPLA_INST_0_68275 : AO1A
      port map(A => HIEFFPLA_NET_0_72704, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, C => 
        HIEFFPLA_NET_0_72691, Y => HIEFFPLA_NET_0_72692);
    
    HIEFFPLA_INST_0_62693 : NOR3A
      port map(A => HIEFFPLA_NET_0_73887, B => 
        HIEFFPLA_NET_0_73909, C => HIEFFPLA_NET_0_73914, Y => 
        HIEFFPLA_NET_0_73927);
    
    HIEFFPLA_INST_0_65277 : AND3C
      port map(A => \Science_0/ADC_READ_0/state[1]_net_1\, B => 
        \Science_0/ADC_READ_0/state[0]_net_1\, C => 
        \Science_0/ADC_READ_0/countere\, Y => 
        HIEFFPLA_NET_0_73426);
    
    \General_Controller_0/constant_bias_voltage_0[11]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[11]_net_1\);
    
    HIEFFPLA_INST_0_66849 : AO1
      port map(A => HIEFFPLA_NET_0_73015, B => 
        HIEFFPLA_NET_0_73097, C => HIEFFPLA_NET_0_73013, Y => 
        HIEFFPLA_NET_0_73022);
    
    \Science_0/ADC_READ_0/exp_packet_1[37]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[3]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[37]\);
    
    HIEFFPLA_INST_0_69667 : OA1A
      port map(A => HIEFFPLA_NET_0_72382, B => 
        \Sensors_0/Pressure_Sensor_0/state[8]\, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_we\, 
        Y => HIEFFPLA_NET_0_72333);
    
    HIEFFPLA_INST_0_62537 : AO1B
      port map(A => HIEFFPLA_NET_0_73974, B => 
        HIEFFPLA_NET_0_73905, C => HIEFFPLA_NET_0_73961, Y => 
        HIEFFPLA_NET_0_73962);
    
    HIEFFPLA_INST_0_69574 : NAND3C
      port map(A => HIEFFPLA_NET_0_72360, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72361);
    
    HIEFFPLA_INST_0_56530 : AX1C
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[1]_net_1\, B
         => 
        \Data_Saving_0/Interrupt_Generator_0/counter[0]_net_1\, C
         => 
        \Data_Saving_0/Interrupt_Generator_0/counter[2]_net_1\, Y
         => HIEFFPLA_NET_0_75251);
    
    HIEFFPLA_INST_0_68896 : AND2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/isSetup_net_1\, B
         => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72528);
    
    \General_Controller_0/sweep_table_samples_per_point[8]\ : 
        DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[8]_net_1\);
    
    HIEFFPLA_INST_0_57252 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[59]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_75111);
    
    HIEFFPLA_INST_0_69867 : NOR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72286);
    
    HIEFFPLA_INST_0_68727 : NAND2B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\, B
         => \Sensors_0/Gyro_0/I2C_Master_0/next_state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72577);
    
    HIEFFPLA_INST_0_68442 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[2]_net_1\, B => 
        HIEFFPLA_NET_0_72646, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, Y => 
        HIEFFPLA_NET_0_72649);
    
    HIEFFPLA_INST_0_66700 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_73060);
    
    HIEFFPLA_INST_0_67408 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, Y
         => HIEFFPLA_NET_0_72889);
    
    \General_Controller_0/status_bits_1[38]\ : DFN1E1
      port map(D => General_Controller_0_en_data_saving, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74266, Q => 
        \Data_Hub_Packets_0_status_packet[5]\);
    
    HIEFFPLA_INST_0_67248 : NAND3C
      port map(A => HIEFFPLA_NET_0_72909, B => 
        HIEFFPLA_NET_0_72770, C => HIEFFPLA_NET_0_72886, Y => 
        HIEFFPLA_NET_0_72928);
    
    HIEFFPLA_INST_0_58668 : AND2
      port map(A => \General_Controller_0_gs_id[7]\, B => 
        HIEFFPLA_NET_0_74484, Y => HIEFFPLA_NET_0_74708);
    
    \Science_0/ADC_READ_0/chan3_data[3]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[3]\);
    
    HIEFFPLA_INST_0_61593 : NAND3C
      port map(A => HIEFFPLA_NET_0_74179, B => 
        HIEFFPLA_NET_0_74178, C => HIEFFPLA_NET_0_73979, Y => 
        HIEFFPLA_NET_0_74177);
    
    HIEFFPLA_INST_0_66492 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73108);
    
    \Communications_0/UART_0/tx_byte[7]\ : DFN1E1
      port map(D => \GS_Readout_0_send[7]\, CLK => CLKINT_0_Y_0, 
        E => HIEFFPLA_NET_0_75504, Q => 
        \Communications_0/UART_0/tx_byte[7]_net_1\);
    
    HIEFFPLA_INST_0_69944 : AO1D
      port map(A => HIEFFPLA_NET_0_72256, B => 
        HIEFFPLA_NET_0_72304, C => HIEFFPLA_NET_0_72251, Y => 
        HIEFFPLA_NET_0_72262);
    
    HIEFFPLA_INST_0_61848 : NOR3B
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        HIEFFPLA_NET_0_73948, C => 
        \General_Controller_0/uc_rx_byte[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74117);
    
    HIEFFPLA_INST_0_61548 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[61]\, B => 
        \Timekeeper_0_milliseconds[21]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74185);
    
    HIEFFPLA_INST_0_54941 : AOI1B
      port map(A => HIEFFPLA_NET_0_75635, B => 
        HIEFFPLA_NET_0_75636, C => HIEFFPLA_NET_0_75631, Y => 
        HIEFFPLA_NET_0_75633);
    
    \General_Controller_0/ext_rx_state[1]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_74299, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \General_Controller_0/ext_rx_state_i_0[1]\);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/data_out_rdy\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72341, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72393, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\);
    
    HIEFFPLA_INST_0_56280 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[10]\\\\\, B
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[9]\\\\\, C
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[8]\\\\\, Y
         => HIEFFPLA_NET_0_75321);
    
    HIEFFPLA_INST_0_55834 : AND2
      port map(A => \Communications_0/UART_1/tx_clk_count_i_0[2]\, 
        B => \Communications_0/UART_1/tx_clk_count_i_0[3]\, Y => 
        HIEFFPLA_NET_0_75416);
    
    HIEFFPLA_INST_0_65775 : XA1B
      port map(A => HIEFFPLA_NET_0_73281, B => 
        \Science_0/ADC_READ_0/cnt[7]_net_1\, C => 
        HIEFFPLA_NET_0_73241, Y => HIEFFPLA_NET_0_73282);
    
    HIEFFPLA_INST_0_63650 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[11]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_samples_per_point[11]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73734);
    
    HIEFFPLA_INST_0_63446 : MX2
      port map(A => HIEFFPLA_NET_0_73754, B => 
        HIEFFPLA_NET_0_73687, S => HIEFFPLA_NET_0_73608, Y => 
        HIEFFPLA_NET_0_73762);
    
    HIEFFPLA_INST_0_57913 : AO1
      port map(A => \Science_0_exp_packet_0[66]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75132, Y => HIEFFPLA_NET_0_74907);
    
    HIEFFPLA_INST_0_55692 : MX2A
      port map(A => HIEFFPLA_NET_0_75445, B => 
        HIEFFPLA_NET_0_75439, S => 
        \Communications_0/UART_1/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75446);
    
    HIEFFPLA_INST_0_55176 : AND2B
      port map(A => \Communications_0/UART_0/rx_clk_count_c0\, B
         => HIEFFPLA_NET_0_75567, Y => HIEFFPLA_NET_0_75568);
    
    \General_Controller_0/command[2]\ : DFN1E1
      port map(D => \Communications_0_ext_recv[2]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74300, Q => 
        \General_Controller_0/command[2]_net_1\);
    
    HIEFFPLA_INST_0_57737 : AO1B
      port map(A => \Sensors_0_acc_time[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74956, Y => HIEFFPLA_NET_0_74957);
    
    HIEFFPLA_INST_0_63166 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state_0[3]_net_1\, 
        B => HIEFFPLA_NET_0_73988, C => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73817);
    
    HIEFFPLA_INST_0_56027 : AND2A
      port map(A => \Data_Saving_0/FPGA_Buffer_0/empty\, B => 
        FMC_NOE_c, Y => \Data_Saving_0/FPGA_Buffer_0/MEMRENEG\);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/temp[6]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72907, Q => 
        \Sensors_0_acc_temp[6]\);
    
    HIEFFPLA_INST_0_65248 : AND3B
      port map(A => \Sensors_0_pressure_raw[22]\, B => 
        \Sensors_0_pressure_raw[20]\, C => HIEFFPLA_NET_0_73428, 
        Y => HIEFFPLA_NET_0_73435);
    
    \General_Controller_0/led1\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74273, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => LED1_c);
    
    HIEFFPLA_INST_0_64648 : AOI1A
      port map(A => HIEFFPLA_NET_0_73612, B => 
        \General_Controller_0/uc_tx_state[7]_net_1\, C => 
        HIEFFPLA_NET_0_73576, Y => HIEFFPLA_NET_0_73577);
    
    HIEFFPLA_INST_0_59175 : AO1C
      port map(A => HIEFFPLA_NET_0_74636, B => 
        HIEFFPLA_NET_0_74580, C => Communications_0_ext_tx_rdy, Y
         => HIEFFPLA_NET_0_74595);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRY[7]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75313, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[7]\\\\\);
    
    HIEFFPLA_INST_0_67746 : NAND3C
      port map(A => HIEFFPLA_NET_0_72730, B => 
        HIEFFPLA_NET_0_72733, C => HIEFFPLA_NET_0_72806, Y => 
        HIEFFPLA_NET_0_72810);
    
    HIEFFPLA_INST_0_69578 : OR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]_net_1\, 
        B => \Sensors_0/Pressure_Sensor_0/state[8]\, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72360);
    
    HIEFFPLA_INST_0_71206 : AND3B
      port map(A => HIEFFPLA_NET_0_71974, B => 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\, C => 
        \Communications_0/UART_1/rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75439);
    
    HIEFFPLA_INST_0_68856 : AOI1
      port map(A => HIEFFPLA_NET_0_72531, B => 
        HIEFFPLA_NET_0_72486, C => HIEFFPLA_NET_0_72522, Y => 
        HIEFFPLA_NET_0_72538);
    
    HIEFFPLA_INST_0_55878 : XO1A
      port map(A => HIEFFPLA_NET_0_75412, B => 
        \Communications_0/UART_1/tx_clk_count_i_0[5]\, C => 
        HIEFFPLA_NET_0_75419, Y => HIEFFPLA_NET_0_75406);
    
    HIEFFPLA_INST_0_66670 : OA1C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        B => HIEFFPLA_NET_0_73144, C => HIEFFPLA_NET_0_73068, Y
         => HIEFFPLA_NET_0_73069);
    
    HIEFFPLA_INST_0_70417 : AX1C
      port map(A => \Timekeeper_0_microseconds[19]\, B => 
        HIEFFPLA_NET_0_72158, C => 
        \Timekeeper_0_microseconds[20]\, Y => 
        HIEFFPLA_NET_0_72139);
    
    HIEFFPLA_INST_0_59225 : NOR3B
      port map(A => \GS_Readout_0/state[4]_net_1\, B => 
        HIEFFPLA_NET_0_74382, C => Communications_0_ext_tx_rdy, Y
         => HIEFFPLA_NET_0_74585);
    
    HIEFFPLA_INST_0_68573 : AOI1C
      port map(A => HIEFFPLA_NET_0_72603, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, Y => 
        HIEFFPLA_NET_0_72614);
    
    HIEFFPLA_INST_0_59039 : NOR3A
      port map(A => HIEFFPLA_NET_0_74662, B => 
        \GS_Readout_0/state[6]_net_1\, C => HIEFFPLA_NET_0_74640, 
        Y => HIEFFPLA_NET_0_74629);
    
    HIEFFPLA_INST_0_66325 : AOI1C
      port map(A => HIEFFPLA_NET_0_73149, B => 
        HIEFFPLA_NET_0_73147, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73145);
    
    HIEFFPLA_INST_0_64297 : MX2
      port map(A => HIEFFPLA_NET_0_73728, B => 
        HIEFFPLA_NET_0_73720, S => HIEFFPLA_NET_0_73619, Y => 
        HIEFFPLA_NET_0_73640);
    
    HIEFFPLA_INST_0_69038 : NOR3A
      port map(A => HIEFFPLA_NET_0_72495, B => 
        HIEFFPLA_NET_0_72548, C => HIEFFPLA_NET_0_72481, Y => 
        HIEFFPLA_NET_0_72489);
    
    HIEFFPLA_INST_0_63746 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[3]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[3]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73718);
    
    HIEFFPLA_INST_0_60935 : OR3A
      port map(A => HIEFFPLA_NET_0_74337, B => 
        \General_Controller_0/flight_state[2]_net_1\, C => 
        \General_Controller_0/flight_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74316);
    
    HIEFFPLA_INST_0_57661 : AO1B
      port map(A => \Sensors_0_gyro_y[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74977, Y => HIEFFPLA_NET_0_74978);
    
    HIEFFPLA_INST_0_60294 : NOR3A
      port map(A => HIEFFPLA_NET_0_74450, B => 
        HIEFFPLA_NET_0_74490, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74435);
    
    HIEFFPLA_INST_0_57830 : AOI1
      port map(A => \Sensors_0_acc_time[18]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74931, Y => HIEFFPLA_NET_0_74932);
    
    \General_Controller_0/constant_bias_voltage_0[13]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[13]_net_1\);
    
    \General_Controller_0/command[4]\ : DFN1E1
      port map(D => \Communications_0_ext_recv[4]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74300, Q => 
        \General_Controller_0/command[4]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/temp[2]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72555, Q => 
        \Sensors_0_gyro_temp[2]\);
    
    HIEFFPLA_INST_0_55955 : NOR2A
      port map(A => HIEFFPLA_NET_0_75381, B => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_75385);
    
    HIEFFPLA_INST_0_59148 : NAND3C
      port map(A => HIEFFPLA_NET_0_74584, B => 
        HIEFFPLA_NET_0_74590, C => HIEFFPLA_NET_0_74616, Y => 
        HIEFFPLA_NET_0_74600);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[0]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72808, Q => 
        \Sensors_0_mag_z[0]\);
    
    HIEFFPLA_INST_0_65467 : AX1
      port map(A => HIEFFPLA_NET_0_73379, B => 
        \Science_0/ADC_READ_0/cnt2dn[5]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt2dn[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73369);
    
    \Data_Saving_0/Interrupt_Generator_0/uC_interrupt\ : DFN1E0C1
      port map(D => 
        \Data_Saving_0/Interrupt_Generator_0/counter[9]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75242, Q => FPGA_BUF_INT_c);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72471, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\);
    
    HIEFFPLA_INST_0_57634 : AOI1
      port map(A => \Science_0_exp_packet_0[32]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74985, Y => HIEFFPLA_NET_0_74986);
    
    HIEFFPLA_INST_0_65746 : XA1B
      port map(A => \Science_0/ADC_READ_0/cnt[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_73241, Y => HIEFFPLA_NET_0_73291);
    
    HIEFFPLA_INST_0_64081 : MX2
      port map(A => HIEFFPLA_NET_0_73636, B => 
        HIEFFPLA_NET_0_73628, S => HIEFFPLA_NET_0_73585, Y => 
        HIEFFPLA_NET_0_73673);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[14]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[14]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[14]\);
    
    HIEFFPLA_INST_0_71015 : AXOI3
      port map(A => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, B => 
        \General_Controller_0/uc_tx_substate[2]_net_1\, C => 
        Communications_0_uc_tx_rdy, Y => HIEFFPLA_NET_0_71988);
    
    HIEFFPLA_INST_0_57350 : AO1A
      port map(A => HIEFFPLA_NET_0_75117, B => 
        \Sensors_0_acc_temp[5]\, C => HIEFFPLA_NET_0_75068, Y => 
        HIEFFPLA_NET_0_75069);
    
    HIEFFPLA_INST_0_64652 : AO1A
      port map(A => HIEFFPLA_NET_0_73605, B => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, C => 
        \General_Controller_0/uc_tx_state[15]_net_1\, Y => 
        HIEFFPLA_NET_0_73576);
    
    HIEFFPLA_INST_0_62159 : AND3C
      port map(A => \General_Controller_0/uc_rx_state_0[1]_net_1\, 
        B => HIEFFPLA_NET_0_73897, C => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74040);
    
    HIEFFPLA_INST_0_56033 : AND3
      port map(A => HIEFFPLA_NET_0_75327, B => 
        HIEFFPLA_NET_0_75360, C => HIEFFPLA_NET_0_75363, Y => 
        HIEFFPLA_NET_0_75364);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1E1C0_data_out[5]\\\\/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75282, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \FMC_DA_c[5]\);
    
    HIEFFPLA_INST_0_62672 : NOR3B
      port map(A => HIEFFPLA_NET_0_74018, B => 
        HIEFFPLA_NET_0_73887, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73931);
    
    HIEFFPLA_INST_0_55538 : NOR2A
      port map(A => \Communications_0/UART_1/rx_count[2]_net_1\, 
        B => \Communications_0/UART_1/rx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75484);
    
    HIEFFPLA_INST_0_59487 : MX2
      port map(A => HIEFFPLA_NET_0_74522, B => 
        HIEFFPLA_NET_0_74572, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74547);
    
    \Eject_Signal_Debounce_0/ms_cnt[1]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74746, CLK => CLKINT_0_Y_0, Q
         => \Eject_Signal_Debounce_0/ms_cnt[1]_net_1\);
    
    HIEFFPLA_INST_0_62798 : AND2
      port map(A => \General_Controller_0/uc_rx_state[4]_net_1\, 
        B => \General_Controller_0/uc_rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73900);
    
    \Science_0/ADC_READ_0/chan1_data[2]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[2]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[7]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72804, Q => 
        \Sensors_0_mag_x[7]\);
    
    HIEFFPLA_INST_0_59875 : MX2
      port map(A => HIEFFPLA_NET_0_74519, B => 
        HIEFFPLA_NET_0_74514, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74493);
    
    HIEFFPLA_INST_0_61081 : NAND3C
      port map(A => \Timekeeper_0_milliseconds[1]\, B => 
        \Timekeeper_0_milliseconds[0]\, C => 
        \Timekeeper_0_milliseconds[2]\, Y => HIEFFPLA_NET_0_74282);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/i2c_addr_1[3]\ : 
        DFN1E0
      port map(D => HIEFFPLA_NET_0_72988, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72774, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[3]\);
    
    HIEFFPLA_INST_0_56456 : XNOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[7]\\\\\, B => 
        HIEFFPLA_NET_0_75321, Y => HIEFFPLA_NET_0_75277);
    
    HIEFFPLA_INST_0_67866 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72784);
    
    HIEFFPLA_INST_0_66854 : AO1
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_73021);
    
    HIEFFPLA_INST_0_58013 : AO1
      port map(A => \Science_0_exp_packet_0[72]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75121, Y => HIEFFPLA_NET_0_74879);
    
    HIEFFPLA_INST_0_55314 : MX2
      port map(A => HIEFFPLA_NET_0_75538, B => 
        HIEFFPLA_NET_0_75537, S => 
        \Communications_0/UART_0/tx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75541);
    
    HIEFFPLA_INST_0_63301 : AO1
      port map(A => HIEFFPLA_NET_0_73810, B => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, C => 
        HIEFFPLA_NET_0_73804, Y => HIEFFPLA_NET_0_73783);
    
    HIEFFPLA_INST_0_61793 : AX1C
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[7]_net_1\, B
         => HIEFFPLA_NET_0_74145, C => 
        \General_Controller_0/sweep_table_sweep_cnt[8]_net_1\, Y
         => HIEFFPLA_NET_0_74130);
    
    \Data_Saving_0/Packet_Saver_0/data_out[17]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75228, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[17]\);
    
    HIEFFPLA_INST_0_63626 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[15]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_sample_skip[15]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73738);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_WADDR[7]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75304, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[7]\\\\\);
    
    HIEFFPLA_INST_0_62797 : NOR2A
      port map(A => \General_Controller_0/uc_rx_state[1]_net_1\, 
        B => \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73901);
    
    HIEFFPLA_INST_0_67664 : AO1E
      port map(A => HIEFFPLA_NET_0_72888, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        C => HIEFFPLA_NET_0_72829, Y => HIEFFPLA_NET_0_72830);
    
    \Data_Saving_0/Packet_Saver_0/packet_select[9]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74775, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[9]\);
    
    HIEFFPLA_INST_0_63818 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[7]_net_1\, 
        B => \General_Controller_0/sweep_table_points[7]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73706);
    
    HIEFFPLA_INST_0_60203 : MX2
      port map(A => HIEFFPLA_NET_0_74470, B => 
        HIEFFPLA_NET_0_74508, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74446);
    
    \LDCS_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => LDCS_c, E => \VCC\, DOUT => 
        \LDCS_pad/U0/NET1\, EOUT => \LDCS_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_62603 : NOR3A
      port map(A => HIEFFPLA_NET_0_73905, B => 
        HIEFFPLA_NET_0_73890, C => HIEFFPLA_NET_0_73781, Y => 
        HIEFFPLA_NET_0_73947);
    
    HIEFFPLA_INST_0_67708 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        B => HIEFFPLA_NET_0_72813, C => HIEFFPLA_NET_0_72752, Y
         => HIEFFPLA_NET_0_72818);
    
    HIEFFPLA_INST_0_56702 : MX2
      port map(A => HIEFFPLA_NET_0_75190, B => 
        HIEFFPLA_NET_0_75050, S => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75223);
    
    HIEFFPLA_INST_0_69896 : NAND3C
      port map(A => HIEFFPLA_NET_0_72278, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72275);
    
    HIEFFPLA_INST_0_58431 : AOI1
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/old_mag_new_data_i_0\, B
         => Sensors_0_mag_new_data, C => 
        \Data_Saving_0/Packet_Saver_0/mag_flag_net_1\, Y => 
        HIEFFPLA_NET_0_74769);
    
    \General_Controller_0/sweep_table_samples_per_step[6]\ : 
        DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[6]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[6]_net_1\);
    
    \Science_0/ADC_READ_0/chan6_data[6]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[6]\);
    
    \Science_0/ADC_READ_0/chan0_data[6]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[6]\);
    
    \General_Controller_0/sweep_table_nof_steps[7]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73980, Q => 
        \General_Controller_0/sweep_table_nof_steps[7]_net_1\);
    
    \General_Controller_0/sweep_table_sweep_cnt[15]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74138, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[15]_net_1\);
    
    HIEFFPLA_INST_0_63936 : MX2
      port map(A => HIEFFPLA_NET_0_73666, B => 
        HIEFFPLA_NET_0_73658, S => HIEFFPLA_NET_0_73594, Y => 
        HIEFFPLA_NET_0_73687);
    
    HIEFFPLA_INST_0_68800 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, B
         => CLKINT_1_Y, C => HIEFFPLA_NET_0_72479, Y => 
        HIEFFPLA_NET_0_72555);
    
    HIEFFPLA_INST_0_69694 : NAND3C
      port map(A => PRESSURE_SCL_c, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[2]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72327);
    
    HIEFFPLA_INST_0_65381 : NOR3B
      port map(A => HIEFFPLA_NET_0_73276, B => 
        HIEFFPLA_NET_0_73393, C => 
        \Science_0/ADC_READ_0/cnt1up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73394);
    
    HIEFFPLA_INST_0_65593 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt3up[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt3up[0]_net_1\, C => 
        HIEFFPLA_NET_0_73338, Y => HIEFFPLA_NET_0_73335);
    
    HIEFFPLA_INST_0_70044 : NAND3
      port map(A => HIEFFPLA_NET_0_72278, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_write_done\, Y
         => HIEFFPLA_NET_0_72236);
    
    HIEFFPLA_INST_0_68286 : NAND2B
      port map(A => HIEFFPLA_NET_0_72690, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_72689);
    
    HIEFFPLA_INST_0_59036 : NAND3C
      port map(A => HIEFFPLA_NET_0_74449, B => 
        HIEFFPLA_NET_0_74628, C => HIEFFPLA_NET_0_74629, Y => 
        HIEFFPLA_NET_0_74630);
    
    \LA0_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => LA0_c, E => \VCC\, DOUT => \LA0_pad/U0/NET1\, 
        EOUT => \LA0_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_59714 : MX2
      port map(A => HIEFFPLA_NET_0_74390, B => 
        HIEFFPLA_NET_0_74427, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74518);
    
    \General_Controller_0/uc_rx_byte[1]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[1]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte[1]_net_1\);
    
    HIEFFPLA_INST_0_62033 : AND2
      port map(A => HIEFFPLA_NET_0_74062, B => 
        HIEFFPLA_NET_0_73956, Y => HIEFFPLA_NET_0_74066);
    
    HIEFFPLA_INST_0_58961 : NAND3C
      port map(A => HIEFFPLA_NET_0_74632, B => 
        HIEFFPLA_NET_0_74639, C => HIEFFPLA_NET_0_74623, Y => 
        HIEFFPLA_NET_0_74648);
    
    HIEFFPLA_INST_0_56487 : AX1C
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\, B
         => HIEFFPLA_NET_0_75257, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[10]\\\\\, Y
         => HIEFFPLA_NET_0_75267);
    
    HIEFFPLA_INST_0_69730 : AND3B
      port map(A => HIEFFPLA_NET_0_72394, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        C => HIEFFPLA_NET_0_72380, Y => HIEFFPLA_NET_0_72320);
    
    HIEFFPLA_INST_0_68989 : AND2
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0_write_done\, B
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        Y => HIEFFPLA_NET_0_72506);
    
    HIEFFPLA_INST_0_56167 : XA1A
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, B
         => HIEFFPLA_NET_0_75370, C => HIEFFPLA_NET_0_75273, Y
         => HIEFFPLA_NET_0_75338);
    
    AFLSDF_INV_13 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_13\);
    
    HIEFFPLA_INST_0_68096 : NOR3B
      port map(A => HIEFFPLA_NET_0_72740, B => 
        HIEFFPLA_NET_0_72929, C => HIEFFPLA_NET_0_72752, Y => 
        HIEFFPLA_NET_0_72730);
    
    HIEFFPLA_INST_0_55619 : XA1
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[25]_net_1\, B => 
        HIEFFPLA_NET_0_75462, C => HIEFFPLA_NET_0_75437, Y => 
        HIEFFPLA_NET_0_75463);
    
    HIEFFPLA_INST_0_57219 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[50]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75123);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[1]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72265, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_65470 : XA1C
      port map(A => \Science_0/ADC_READ_0/cnt2dn[7]_net_1\, B => 
        HIEFFPLA_NET_0_73386, C => HIEFFPLA_NET_0_73381, Y => 
        HIEFFPLA_NET_0_73368);
    
    HIEFFPLA_INST_0_69209 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, B
         => HIEFFPLA_NET_0_72445, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        Y => HIEFFPLA_NET_0_72446);
    
    \Science_0/ADC_READ_0/chan4_data[8]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[8]\);
    
    HIEFFPLA_INST_0_69850 : AO1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        B => HIEFFPLA_NET_0_72244, C => HIEFFPLA_NET_0_72289, Y
         => HIEFFPLA_NET_0_72291);
    
    HIEFFPLA_INST_0_67055 : NAND2B
      port map(A => \Sensors_0/Accelerometer_0/state_0[8]\, B => 
        HIEFFPLA_NET_0_72735, Y => HIEFFPLA_NET_0_72977);
    
    HIEFFPLA_INST_0_62401 : NAND3C
      port map(A => HIEFFPLA_NET_0_73989, B => 
        HIEFFPLA_NET_0_74099, C => HIEFFPLA_NET_0_73889, Y => 
        HIEFFPLA_NET_0_73990);
    
    HIEFFPLA_INST_0_68925 : OA1A
      port map(A => HIEFFPLA_NET_0_72518, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/isSetup_net_1\, C
         => HIEFFPLA_NET_0_72519, Y => HIEFFPLA_NET_0_72520);
    
    HIEFFPLA_INST_0_66818 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_73025, C => ACCE_SCL_c, Y => 
        HIEFFPLA_NET_0_73028);
    
    HIEFFPLA_INST_0_58819 : NOR3B
      port map(A => HIEFFPLA_NET_0_74433, B => 
        HIEFFPLA_NET_0_74633, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74680);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[5]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[5]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[5]\);
    
    \Pressure_Signal_Debounce_0/ms_cnt[2]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73493, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[2]_net_1\);
    
    HIEFFPLA_INST_0_69887 : AND3
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72279);
    
    HIEFFPLA_INST_0_70943 : OA1C
      port map(A => HIEFFPLA_NET_0_72003, B => 
        HIEFFPLA_NET_0_72761, C => HIEFFPLA_NET_0_72933, Y => 
        HIEFFPLA_NET_0_72978);
    
    \Communications_0/UART_0/rx_count[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75559, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75555, Q => 
        \Communications_0/UART_0/rx_count[2]_net_1\);
    
    HIEFFPLA_INST_0_57947 : AO1B
      port map(A => \Sensors_0_mag_time[14]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74896, Y => HIEFFPLA_NET_0_74897);
    
    \General_Controller_0/constant_bias_voltage_0[14]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[14]_net_1\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73029, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\);
    
    \General_Controller_0/constant_bias_voltage_0[12]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[12]_net_1\);
    
    HIEFFPLA_INST_0_69993 : NOR3B
      port map(A => HIEFFPLA_NET_0_72238, B => 
        HIEFFPLA_NET_0_72285, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72250);
    
    HIEFFPLA_INST_0_67961 : NOR3A
      port map(A => HIEFFPLA_NET_0_72881, B => 
        HIEFFPLA_NET_0_72739, C => HIEFFPLA_NET_0_72888, Y => 
        HIEFFPLA_NET_0_72766);
    
    \Science_0/ADC_READ_0/data_b[13]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[13]_net_1\);
    
    HIEFFPLA_INST_0_62811 : NAND2B
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73897);
    
    HIEFFPLA_INST_0_67137 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[6]_net_1\, 
        Y => HIEFFPLA_NET_0_72956);
    
    HIEFFPLA_INST_0_64667 : AND2
      port map(A => 
        \General_Controller_0/uc_tx_nextstate[1]_net_1\, B => 
        HIEFFPLA_NET_0_73584, Y => HIEFFPLA_NET_0_73572);
    
    HIEFFPLA_INST_0_68918 : OA1A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, B
         => \Sensors_0/Gyro_0/I2C_Master_0_s_ack_error\, C => 
        HIEFFPLA_NET_0_72516, Y => HIEFFPLA_NET_0_72522);
    
    HIEFFPLA_INST_0_56483 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[5]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[4]\\\\\, Y => 
        HIEFFPLA_NET_0_75269);
    
    \General_Controller_0/gs_id[4]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73922, Q => 
        \General_Controller_0_gs_id[4]\);
    
    HIEFFPLA_INST_0_61866 : NOR3B
      port map(A => HIEFFPLA_NET_0_74094, B => 
        \General_Controller_0/uc_rx_state[0]_net_1\, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74113);
    
    HIEFFPLA_INST_0_56952 : MX2
      port map(A => HIEFFPLA_NET_0_74972, B => 
        HIEFFPLA_NET_0_74903, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75191);
    
    HIEFFPLA_INST_0_57287 : AND2
      port map(A => \Sensors_0_acc_time[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, Y
         => HIEFFPLA_NET_0_75093);
    
    HIEFFPLA_INST_0_57505 : AO1
      port map(A => \Sensors_0_acc_z[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74837, Y => HIEFFPLA_NET_0_75026);
    
    \General_Controller_0/command[0]\ : DFN1E1
      port map(D => \Communications_0_ext_recv[0]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74300, Q => 
        \General_Controller_0/command[0]_net_1\);
    
    HIEFFPLA_INST_0_66279 : NAND2
      port map(A => HIEFFPLA_NET_0_73179, B => 
        \Science_0/SET_LP_GAIN_0/state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73158);
    
    \General_Controller_0/sweep_table_sweep_cnt[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74135, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[3]_net_1\);
    
    AFLSDF_INV_16 : INV
      port map(A => Sensors_0_gyro_new_data, Y => \AFLSDF_INV_16\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[4]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[4]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[4]\);
    
    HIEFFPLA_INST_0_58581 : AX1C
      port map(A => HIEFFPLA_NET_0_74729, B => 
        \Eject_Signal_Debounce_0/ms_cnt[1]_net_1\, C => 
        \Eject_Signal_Debounce_0/ms_cnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74730);
    
    HIEFFPLA_INST_0_57716 : AOI1
      port map(A => \Science_0_exp_packet_0[56]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74822, Y => HIEFFPLA_NET_0_74961);
    
    HIEFFPLA_INST_0_57135 : AND2
      port map(A => \Sensors_0_acc_y[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        Y => HIEFFPLA_NET_0_75162);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]\ : 
        DFN1P1
      port map(D => HIEFFPLA_NET_0_72746, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\);
    
    HIEFFPLA_INST_0_56386 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[1]\\\\\, B
         => HIEFFPLA_NET_0_75293, Y => HIEFFPLA_NET_0_75294);
    
    HIEFFPLA_INST_0_69521 : MX2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[1]\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[3]\, 
        S => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72372);
    
    HIEFFPLA_INST_0_68121 : MX2
      port map(A => HIEFFPLA_NET_0_72723, B => 
        HIEFFPLA_NET_0_72713, S => HIEFFPLA_NET_0_72876, Y => 
        HIEFFPLA_NET_0_72727);
    
    HIEFFPLA_INST_0_67787 : XO1A
      port map(A => HIEFFPLA_NET_0_72737, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72802);
    
    HIEFFPLA_INST_0_67843 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72789);
    
    HIEFFPLA_INST_0_67672 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, B
         => HIEFFPLA_NET_0_72734, C => HIEFFPLA_NET_0_72743, Y
         => HIEFFPLA_NET_0_72827);
    
    HIEFFPLA_INST_0_63325 : NAND3C
      port map(A => HIEFFPLA_NET_0_73811, B => 
        HIEFFPLA_NET_0_73804, C => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73776);
    
    HIEFFPLA_INST_0_61884 : NAND3
      port map(A => HIEFFPLA_NET_0_74074, B => 
        HIEFFPLA_NET_0_74081, C => 
        \General_Controller_0/uc_rx_byte[7]_net_1\, Y => 
        HIEFFPLA_NET_0_74109);
    
    \I2C_PassThrough_0/cnt[4]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73516, CLK => CLKINT_0_Y_0, Q
         => \I2C_PassThrough_0/cnt[4]_net_1\);
    
    HIEFFPLA_INST_0_69032 : NOR3A
      port map(A => HIEFFPLA_NET_0_72496, B => 
        HIEFFPLA_NET_0_72548, C => HIEFFPLA_NET_0_72481, Y => 
        HIEFFPLA_NET_0_72490);
    
    HIEFFPLA_INST_0_68839 : AO1
      port map(A => General_Controller_0_en_sensors, B => 
        \Sensors_0/Gyro_0/state[8]\, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, Y
         => HIEFFPLA_NET_0_72543);
    
    HIEFFPLA_INST_0_66822 : NOR3A
      port map(A => HIEFFPLA_NET_0_73144, B => 
        HIEFFPLA_NET_0_73060, C => ACCE_SCL_c, Y => 
        HIEFFPLA_NET_0_73027);
    
    HIEFFPLA_INST_0_63978 : MX2
      port map(A => HIEFFPLA_NET_0_73654, B => 
        HIEFFPLA_NET_0_73646, S => HIEFFPLA_NET_0_73599, Y => 
        HIEFFPLA_NET_0_73683);
    
    HIEFFPLA_INST_0_61444 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[48]\, B => 
        \Timekeeper_0_milliseconds[8]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74198);
    
    AFLSDF_INV_25 : INV
      port map(A => \s_clks_net_0[24]\, Y => \AFLSDF_INV_25\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[8]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75259, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[0]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72783, Q => 
        \Sensors_0_mag_y[0]\);
    
    HIEFFPLA_INST_0_70989 : AXOI2
      port map(A => HIEFFPLA_NET_0_73258, B => 
        HIEFFPLA_NET_0_73382, C => \Science_0/ADC_READ_0_G2[1]\, 
        Y => HIEFFPLA_NET_0_71995);
    
    HIEFFPLA_INST_0_67798 : OR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72799);
    
    HIEFFPLA_INST_0_68268 : NAND3C
      port map(A => HIEFFPLA_NET_0_72625, B => 
        HIEFFPLA_NET_0_72692, C => HIEFFPLA_NET_0_72671, Y => 
        HIEFFPLA_NET_0_72693);
    
    HIEFFPLA_INST_0_59409 : MX2
      port map(A => \Science_0_chan7_data[11]\, B => 
        \Science_0_chan6_data[3]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74558);
    
    HIEFFPLA_INST_0_69130 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[5]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[6]_net_1\, 
        C => HIEFFPLA_NET_0_72557, Y => HIEFFPLA_NET_0_72464);
    
    HIEFFPLA_INST_0_57960 : AOI1
      port map(A => \Sensors_0_gyro_time[15]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74892, Y => HIEFFPLA_NET_0_74893);
    
    \General_Controller_0/sweep_table_write_value[6]\ : DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[6]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[6]_net_1\);
    
    HIEFFPLA_INST_0_69091 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[1]_net_1\, 
        C => HIEFFPLA_NET_0_72556, Y => HIEFFPLA_NET_0_72472);
    
    HIEFFPLA_INST_0_66687 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]_net_1\, 
        B => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73064);
    
    HIEFFPLA_INST_0_57297 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[47]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75086);
    
    \General_Controller_0/st_raddr[4]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[4]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73979, Q => 
        \General_Controller_0_st_raddr_1[4]\);
    
    HIEFFPLA_INST_0_65294 : NOR3B
      port map(A => \Science_0/ADC_READ_0/newflag_net_1\, B => 
        \Science_0/ADC_READ_0/chan[0]_net_1\, C => 
        \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73420);
    
    HIEFFPLA_INST_0_71432 : AX1E
      port map(A => \Science_0/ADC_READ_0/cnt2up[4]_net_1\, B => 
        HIEFFPLA_NET_0_73276, C => \Science_0/ADC_READ_0_G2[0]\, 
        Y => HIEFFPLA_NET_0_71968);
    
    HIEFFPLA_INST_0_69601 : NOR3A
      port map(A => HIEFFPLA_NET_0_72430, B => CLKINT_1_Y, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72353);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/data_out[1]\ : 
        DFN0E1C1
      port map(D => ACCE_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73124, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\);
    
    HIEFFPLA_INST_0_60678 : XA1
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, C => 
        HIEFFPLA_NET_0_74575, Y => HIEFFPLA_NET_0_74378);
    
    HIEFFPLA_INST_0_55936 : AO1A
      port map(A => HIEFFPLA_NET_0_75420, B => 
        HIEFFPLA_NET_0_75394, C => HIEFFPLA_NET_0_75390, Y => 
        HIEFFPLA_NET_0_75391);
    
    HIEFFPLA_INST_0_63161 : OR3B
      port map(A => HIEFFPLA_NET_0_74113, B => 
        HIEFFPLA_NET_0_74074, C => 
        \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73818);
    
    \CLOCK_pad/U0/U1\ : IOIN_IB
      port map(YIN => \CLOCK_pad/U0/NET1\, Y => CLOCK_c);
    
    \Science_0/ADC_READ_0/exp_packet_1[79]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[23]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[79]\);
    
    HIEFFPLA_INST_0_62017 : OR2A
      port map(A => 
        \General_Controller_0/uc_rx_prev_state[4]_net_1\, B => 
        Communications_0_uc_rx_rdy, Y => HIEFFPLA_NET_0_74071);
    
    HIEFFPLA_INST_0_61758 : AND3
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[5]_net_1\, B
         => HIEFFPLA_NET_0_74150, C => 
        \General_Controller_0/sweep_table_sweep_cnt[6]_net_1\, Y
         => HIEFFPLA_NET_0_74145);
    
    \Science_0/ADC_READ_0/chan7_data[6]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[6]\);
    
    \General_Controller_0/status_bits_1[51]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74195, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[51]\);
    
    HIEFFPLA_INST_0_64964 : AND3
      port map(A => \I2C_PassThrough_0/cnt[1]_net_1\, B => 
        \I2C_PassThrough_0/cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_73514, Y => HIEFFPLA_NET_0_73501);
    
    \GS_Readout_0/send[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74710, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74630, Q => 
        \GS_Readout_0_send[6]\);
    
    \General_Controller_0/uc_tx_state[5]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73568, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[5]_net_1\);
    
    HIEFFPLA_INST_0_70421 : AX1C
      port map(A => HIEFFPLA_NET_0_72160, B => 
        \Timekeeper_0_microseconds[21]\, C => 
        \Timekeeper_0_microseconds[22]\, Y => 
        HIEFFPLA_NET_0_72137);
    
    HIEFFPLA_INST_0_70236 : AND3C
      port map(A => HIEFFPLA_NET_0_72311, B => 
        HIEFFPLA_NET_0_72308, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72189);
    
    HIEFFPLA_INST_0_64876 : AND3B
      port map(A => HIEFFPLA_NET_0_73523, B => 
        HIEFFPLA_NET_0_73526, C => HIEFFPLA_NET_0_73528, Y => 
        HIEFFPLA_NET_0_73520);
    
    \Timing_0/s_time[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72046, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_time[4]_net_1\);
    
    HIEFFPLA_INST_0_62708 : NAND3C
      port map(A => HIEFFPLA_NET_0_73890, B => 
        HIEFFPLA_NET_0_73884, C => HIEFFPLA_NET_0_73776, Y => 
        HIEFFPLA_NET_0_73924);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[2]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[2]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[2]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[8]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[8]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[8]\);
    
    HIEFFPLA_INST_0_61963 : AND3C
      port map(A => HIEFFPLA_NET_0_74001, B => 
        HIEFFPLA_NET_0_74002, C => HIEFFPLA_NET_0_74078, Y => 
        HIEFFPLA_NET_0_74088);
    
    \General_Controller_0/gs_id[7]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73922, Q => 
        \General_Controller_0_gs_id[7]\);
    
    HIEFFPLA_INST_0_62745 : AND3A
      port map(A => HIEFFPLA_NET_0_73875, B => 
        \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        \General_Controller_0/uc_rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73915);
    
    HIEFFPLA_INST_0_64972 : AND3
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[5]_net_1\, 
        B => \Pressure_Signal_Debounce_0/ms_cnt[6]_net_1\, C => 
        HIEFFPLA_NET_0_73498, Y => HIEFFPLA_NET_0_73499);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[6]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72800, Q => 
        \Sensors_0_acc_x[6]\);
    
    HIEFFPLA_INST_0_65159 : OA1C
      port map(A => \Sensors_0_pressure_raw[20]\, B => 
        HIEFFPLA_NET_0_73456, C => \Sensors_0_pressure_raw[21]\, 
        Y => HIEFFPLA_NET_0_73455);
    
    \General_Controller_0/sweep_table_samples_per_point[1]\ : 
        DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[1]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[1]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[18]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[18]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[18]\);
    
    HIEFFPLA_INST_0_70486 : AX1C
      port map(A => \Timekeeper_0_milliseconds[9]\, B => 
        HIEFFPLA_NET_0_72124, C => 
        \Timekeeper_0_milliseconds[10]\, Y => 
        HIEFFPLA_NET_0_72115);
    
    \General_Controller_0/constant_bias_voltage_0[3]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[3]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[3]_net_1\);
    
    HIEFFPLA_INST_0_68970 : AO1
      port map(A => HIEFFPLA_NET_0_72509, B => 
        HIEFFPLA_NET_0_72543, C => HIEFFPLA_NET_0_72523, Y => 
        HIEFFPLA_NET_0_72510);
    
    HIEFFPLA_INST_0_69230 : AO1
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]_net_1\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, C => 
        HIEFFPLA_NET_0_72434, Y => HIEFFPLA_NET_0_72443);
    
    HIEFFPLA_INST_0_57585 : AO1B
      port map(A => \Sensors_0_gyro_x[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75000, Y => HIEFFPLA_NET_0_75001);
    
    HIEFFPLA_INST_0_66984 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[2]\, 
        C => HIEFFPLA_NET_0_72884, Y => HIEFFPLA_NET_0_72990);
    
    HIEFFPLA_INST_0_59188 : OR2A
      port map(A => HIEFFPLA_NET_0_74718, B => 
        \GS_Readout_0/prevState[5]_net_1\, Y => 
        HIEFFPLA_NET_0_74592);
    
    HIEFFPLA_INST_0_58482 : AND2
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[1]_net_1\, B => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74754);
    
    HIEFFPLA_INST_0_70247 : NOR3A
      port map(A => HIEFFPLA_NET_0_72185, B => 
        HIEFFPLA_NET_0_72311, C => 
        \Sensors_0/Pressure_Sensor_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72187);
    
    HIEFFPLA_INST_0_60278 : MX2
      port map(A => \Science_0_chan2_data[5]\, B => 
        \Science_0_chan2_data[9]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74438);
    
    HIEFFPLA_INST_0_59173 : NAND3C
      port map(A => HIEFFPLA_NET_0_74360, B => 
        HIEFFPLA_NET_0_74387, C => 
        \GS_Readout_0/subState[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74596);
    
    HIEFFPLA_INST_0_56342 : XOR2
      port map(A => HIEFFPLA_NET_0_75288, B => 
        HIEFFPLA_NET_0_75304, Y => HIEFFPLA_NET_0_75305);
    
    HIEFFPLA_INST_0_57479 : AO1
      port map(A => \Science_0_exp_packet_0[18]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74862, Y => HIEFFPLA_NET_0_75034);
    
    \Science_0/ADC_READ_0/chan3_data[1]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[1]\);
    
    HIEFFPLA_INST_0_66208 : MX2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G1[0]_net_1\, B
         => \Science_0/ADC_READ_0_G1[0]\, S => 
        \Science_0/SET_LP_GAIN_0/state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73177);
    
    \Communications_0/UART_1/recv[0]\ : DFN1E1C1
      port map(D => \Communications_0/UART_1/rx_byte[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75441, Q => \Communications_0_uc_recv[0]\);
    
    \General_Controller_0/sweep_table_points[8]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[8]_net_1\);
    
    HIEFFPLA_INST_0_61961 : AO1E
      port map(A => HIEFFPLA_NET_0_73818, B => 
        HIEFFPLA_NET_0_73819, C => HIEFFPLA_NET_0_74088, Y => 
        HIEFFPLA_NET_0_74089);
    
    HIEFFPLA_INST_0_57693 : AO1
      port map(A => \Sensors_0_pressure_raw[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74848, Y => HIEFFPLA_NET_0_74968);
    
    HIEFFPLA_INST_0_57218 : AND2
      port map(A => \Sensors_0_acc_time[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, Y
         => HIEFFPLA_NET_0_75124);
    
    \General_Controller_0/sweep_table_points[14]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[14]_net_1\);
    
    \Science_0/ADC_READ_0/cnt1dn[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73404, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1dn[4]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[59]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[3]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[59]\);
    
    HIEFFPLA_INST_0_55252 : OA1C
      port map(A => HIEFFPLA_NET_0_75583, B => 
        \Communications_0/UART_0/rx_state[0]_net_1\, C => 
        HIEFFPLA_NET_0_75553, Y => HIEFFPLA_NET_0_75552);
    
    HIEFFPLA_INST_0_62850 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state[1]_net_1\, 
        B => \General_Controller_0/uc_rx_state[0]_net_1\, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73882);
    
    HIEFFPLA_INST_0_61236 : AND2B
      port map(A => HIEFFPLA_NET_0_74217, B => 
        \General_Controller_0/state_seconds[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74240);
    
    HIEFFPLA_INST_0_66038 : XA1B
      port map(A => \Science_0/DAC_SET_0/ADR[0]_net_1\, B => 
        HIEFFPLA_NET_0_73226, C => 
        \Science_0/DAC_SET_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73229);
    
    HIEFFPLA_INST_0_61061 : OR3A
      port map(A => HIEFFPLA_NET_0_74274, B => 
        HIEFFPLA_NET_0_74313, C => HIEFFPLA_NET_0_74283, Y => 
        HIEFFPLA_NET_0_74284);
    
    HIEFFPLA_INST_0_65432 : NAND3
      port map(A => \Science_0/ADC_READ_0/cnt2dn[2]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2dn[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt2dn[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73377);
    
    HIEFFPLA_INST_0_57595 : AO1B
      port map(A => \Sensors_0_acc_x[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74997, Y => HIEFFPLA_NET_0_74998);
    
    \General_Controller_0/sweep_table_probe_id[1]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73924, Q => 
        \General_Controller_0/sweep_table_probe_id[1]_net_1\);
    
    HIEFFPLA_INST_0_62055 : XO1
      port map(A => 
        \General_Controller_0/uc_rx_prev_state[1]_net_1\, B => 
        \General_Controller_0/uc_rx_prev_state[0]_net_1\, C => 
        Communications_0_uc_rx_rdy, Y => HIEFFPLA_NET_0_74062);
    
    HIEFFPLA_INST_0_61939 : OR3A
      port map(A => \General_Controller_0/uc_rx_byte[5]_net_1\, B
         => \General_Controller_0/uc_rx_byte[0]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[6]_net_1\, Y => 
        HIEFFPLA_NET_0_74093);
    
    HIEFFPLA_INST_0_61645 : MX2
      port map(A => \SweepTable_0_RD[12]\, B => 
        \SweepTable_1_RD[12]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74167);
    
    \General_Controller_0/uc_tx_nextstate[0]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73971, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73857, Q => 
        \General_Controller_0/uc_tx_nextstate[0]_net_1\);
    
    HIEFFPLA_INST_0_64973 : AND2
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[9]_net_1\, 
        B => \Pressure_Signal_Debounce_0/ms_cnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73498);
    
    HIEFFPLA_INST_0_58051 : AND2
      port map(A => \Science_0_exp_packet_0[39]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        Y => HIEFFPLA_NET_0_74869);
    
    \General_Controller_0/constant_bias_voltage_0[5]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[5]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[5]_net_1\);
    
    \Communications_0/UART_1/recv[2]\ : DFN1E1C1
      port map(D => \Communications_0/UART_1/rx_byte[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75441, Q => \Communications_0_uc_recv[2]\);
    
    HIEFFPLA_INST_0_67917 : AO1
      port map(A => HIEFFPLA_NET_0_72888, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        C => HIEFFPLA_NET_0_72928, Y => HIEFFPLA_NET_0_72773);
    
    \General_Controller_0/sweep_table_write_value[9]\ : DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[9]_net_1\);
    
    HIEFFPLA_INST_0_62961 : OR2A
      port map(A => HIEFFPLA_NET_0_73938, B => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_73857);
    
    HIEFFPLA_INST_0_65386 : NOR3B
      port map(A => HIEFFPLA_NET_0_73390, B => 
        HIEFFPLA_NET_0_73276, C => 
        \Science_0/ADC_READ_0/cnt1up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73392);
    
    HIEFFPLA_INST_0_70409 : XOR2
      port map(A => HIEFFPLA_NET_0_72162, B => 
        \Timekeeper_0_microseconds[17]\, Y => 
        HIEFFPLA_NET_0_72143);
    
    \General_Controller_0/unit_id[3]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73990, Q => 
        \General_Controller_0_unit_id[3]\);
    
    HIEFFPLA_INST_0_67145 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72953);
    
    HIEFFPLA_INST_0_70770 : OA1A
      port map(A => HIEFFPLA_NET_0_72301, B => 
        HIEFFPLA_NET_0_72235, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72015);
    
    HIEFFPLA_INST_0_60776 : NAND2B
      port map(A => \GS_Readout_0/subState[2]_net_1\, B => 
        \GS_Readout_0/subState[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74360);
    
    HIEFFPLA_INST_0_70575 : AX1C
      port map(A => HIEFFPLA_NET_0_72032, B => 
        \Timing_0/m_count[3]_net_1\, C => 
        \Timing_0/m_count[4]_net_1\, Y => HIEFFPLA_NET_0_72075);
    
    \Science_0/ADC_READ_0/chan1_data[9]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[9]\);
    
    HIEFFPLA_INST_0_56582 : MX2
      port map(A => HIEFFPLA_NET_0_75202, B => 
        HIEFFPLA_NET_0_75077, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75235);
    
    HIEFFPLA_INST_0_57710 : AND3C
      port map(A => HIEFFPLA_NET_0_75153, B => 
        HIEFFPLA_NET_0_74869, C => HIEFFPLA_NET_0_74872, Y => 
        HIEFFPLA_NET_0_74963);
    
    HIEFFPLA_INST_0_66344 : MX2A
      port map(A => HIEFFPLA_NET_0_73135, B => 
        HIEFFPLA_NET_0_73011, S => HIEFFPLA_NET_0_73063, Y => 
        HIEFFPLA_NET_0_73141);
    
    HIEFFPLA_INST_0_55033 : AND3B
      port map(A => HIEFFPLA_NET_0_75562, B => 
        \Communications_0/UART_0/rx_count[2]_net_1\, C => 
        HIEFFPLA_NET_0_75604, Y => HIEFFPLA_NET_0_75609);
    
    HIEFFPLA_INST_0_60258 : MX2
      port map(A => HIEFFPLA_NET_0_74573, B => 
        HIEFFPLA_NET_0_74409, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74440);
    
    HIEFFPLA_INST_0_54985 : XOR2
      port map(A => \General_Controller_0_unit_id[0]\, B => 
        \Communications_0/UART_0_recv[0]\, Y => 
        HIEFFPLA_NET_0_75620);
    
    \General_Controller_0/sweep_table_samples_per_point[10]\ : 
        DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[10]_net_1\);
    
    HIEFFPLA_INST_0_57265 : AND2
      port map(A => \Sensors_0_acc_y[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        Y => HIEFFPLA_NET_0_75104);
    
    HIEFFPLA_INST_0_67905 : OR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72776);
    
    HIEFFPLA_INST_0_67321 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, C
         => CLKINT_1_Y, Y => HIEFFPLA_NET_0_72908);
    
    HIEFFPLA_INST_0_63078 : AND2
      port map(A => \General_Controller_0/uc_rx_byte[3]_net_1\, B
         => \General_Controller_0/uc_rx_byte[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73834);
    
    HIEFFPLA_INST_0_66428 : AND3B
      port map(A => HIEFFPLA_NET_0_73121, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73124);
    
    HIEFFPLA_INST_0_71006 : NAND3C
      port map(A => HIEFFPLA_NET_0_71992, B => 
        HIEFFPLA_NET_0_73480, C => HIEFFPLA_NET_0_73437, Y => 
        HIEFFPLA_NET_0_73479);
    
    HIEFFPLA_INST_0_57114 : NAND3C
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        C => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75165);
    
    HIEFFPLA_INST_0_69677 : AND3
      port map(A => HIEFFPLA_NET_0_72346, B => 
        HIEFFPLA_NET_0_72389, C => HIEFFPLA_NET_0_72410, Y => 
        HIEFFPLA_NET_0_72331);
    
    HIEFFPLA_INST_0_55107 : AND3B
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[25]_net_1\, B => 
        \Communications_0/UART_0/rx_clk_count[26]_net_1\, C => 
        HIEFFPLA_NET_0_75588, Y => HIEFFPLA_NET_0_75589);
    
    HIEFFPLA_INST_0_62191 : NOR3B
      port map(A => HIEFFPLA_NET_0_74018, B => 
        HIEFFPLA_NET_0_73975, C => HIEFFPLA_NET_0_73781, Y => 
        HIEFFPLA_NET_0_74033);
    
    HIEFFPLA_INST_0_59233 : AND3C
      port map(A => HIEFFPLA_NET_0_74382, B => 
        \GS_Readout_0/state[0]_net_1\, C => 
        \GS_Readout_0/state[6]_net_1\, Y => HIEFFPLA_NET_0_74583);
    
    HIEFFPLA_INST_0_56054 : XOR3
      port map(A => HIEFFPLA_NET_0_75269, B => 
        HIEFFPLA_NET_0_75323, C => HIEFFPLA_NET_0_75261, Y => 
        HIEFFPLA_NET_0_75359);
    
    HIEFFPLA_INST_0_55574 : AND3
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[25]_net_1\, B => 
        HIEFFPLA_NET_0_75470, C => 
        \Communications_0/UART_1/rx_clk_count[26]_net_1\, Y => 
        HIEFFPLA_NET_0_75477);
    
    HIEFFPLA_INST_0_64071 : MX2
      port map(A => HIEFFPLA_NET_0_73637, B => 
        HIEFFPLA_NET_0_73629, S => HIEFFPLA_NET_0_73585, Y => 
        HIEFFPLA_NET_0_73674);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_72417, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\);
    
    HIEFFPLA_INST_0_66360 : NAND2
      port map(A => HIEFFPLA_NET_0_73063, B => 
        HIEFFPLA_NET_0_73137, Y => HIEFFPLA_NET_0_73138);
    
    HIEFFPLA_INST_0_69322 : AOI1C
      port map(A => HIEFFPLA_NET_0_72414, B => 
        HIEFFPLA_NET_0_72413, C => HIEFFPLA_NET_0_72355, Y => 
        HIEFFPLA_NET_0_72419);
    
    HIEFFPLA_INST_0_65275 : NAND2B
      port map(A => \Sensors_0_pressure_raw[9]\, B => 
        \Sensors_0_pressure_raw[8]\, Y => HIEFFPLA_NET_0_73427);
    
    \SweepTable_1/SweepTable_R0C0\ : RAM512X18
      port map(RADDR8 => AFLSDF_GND, RADDR7 => 
        \TableSelect_0_RADDR[7]\, RADDR6 => 
        \TableSelect_0_RADDR[6]\, RADDR5 => 
        \TableSelect_0_RADDR[5]\, RADDR4 => 
        \TableSelect_0_RADDR[4]\, RADDR3 => 
        \TableSelect_0_RADDR[3]\, RADDR2 => 
        \TableSelect_0_RADDR[2]\, RADDR1 => 
        \TableSelect_0_RADDR[1]\, RADDR0 => 
        \TableSelect_0_RADDR[0]\, WADDR8 => AFLSDF_GND, WADDR7
         => \General_Controller_0_st_waddr[7]\, WADDR6 => 
        \General_Controller_0_st_waddr[6]\, WADDR5 => 
        \General_Controller_0_st_waddr[5]\, WADDR4 => 
        \General_Controller_0_st_waddr[4]\, WADDR3 => 
        \General_Controller_0_st_waddr[3]\, WADDR2 => 
        \General_Controller_0_st_waddr[2]\, WADDR1 => 
        \General_Controller_0_st_waddr[1]\, WADDR0 => 
        \General_Controller_0_st_waddr[0]\, WD17 => \GND\, WD16
         => \General_Controller_0_st_wdata[15]\, WD15 => 
        \General_Controller_0_st_wdata[14]\, WD14 => 
        \General_Controller_0_st_wdata[13]\, WD13 => 
        \General_Controller_0_st_wdata[12]\, WD12 => 
        \General_Controller_0_st_wdata[11]\, WD11 => 
        \General_Controller_0_st_wdata[10]\, WD10 => 
        \General_Controller_0_st_wdata[9]\, WD9 => 
        \General_Controller_0_st_wdata[8]\, WD8 => \GND\, WD7 => 
        \General_Controller_0_st_wdata[7]\, WD6 => 
        \General_Controller_0_st_wdata[6]\, WD5 => 
        \General_Controller_0_st_wdata[5]\, WD4 => 
        \General_Controller_0_st_wdata[4]\, WD3 => 
        \General_Controller_0_st_wdata[3]\, WD2 => 
        \General_Controller_0_st_wdata[2]\, WD1 => 
        \General_Controller_0_st_wdata[1]\, WD0 => 
        \General_Controller_0_st_wdata[0]\, RW0 => \GND\, RW1 => 
        \VCC\, WW0 => \GND\, WW1 => \VCC\, PIPE => \VCC\, REN => 
        \SweepTable_1.WEBP\, WEN => \SweepTable_1.WEAP\, RCLK => 
        CLKINT_0_Y_0, WCLK => CLKINT_0_Y_0, RESET => 
        \AFLSDF_INV_6\, RD17 => OPEN, RD16 => 
        \SweepTable_1_RD[15]\, RD15 => \SweepTable_1_RD[14]\, 
        RD14 => \SweepTable_1_RD[13]\, RD13 => 
        \SweepTable_1_RD[12]\, RD12 => \SweepTable_1_RD[11]\, 
        RD11 => \SweepTable_1_RD[10]\, RD10 => 
        \SweepTable_1_RD[9]\, RD9 => \SweepTable_1_RD[8]\, RD8
         => OPEN, RD7 => \SweepTable_1_RD[7]\, RD6 => 
        \SweepTable_1_RD[6]\, RD5 => \SweepTable_1_RD[5]\, RD4
         => \SweepTable_1_RD[4]\, RD3 => \SweepTable_1_RD[3]\, 
        RD2 => \SweepTable_1_RD[2]\, RD1 => \SweepTable_1_RD[1]\, 
        RD0 => \SweepTable_1_RD[0]\);
    
    \General_Controller_0/uc_tx_nextstate[5]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73972, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73857, Q => 
        \General_Controller_0/uc_tx_nextstate[5]_net_1\);
    
    HIEFFPLA_INST_0_68639 : XA1A
      port map(A => HIEFFPLA_NET_0_72577, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, C
         => HIEFFPLA_NET_0_72589, Y => HIEFFPLA_NET_0_72599);
    
    HIEFFPLA_INST_0_65145 : AOI1D
      port map(A => \Sensors_0_pressure_raw[9]\, B => 
        \Sensors_0_pressure_raw[8]\, C => 
        \Sensors_0_pressure_raw[11]\, Y => HIEFFPLA_NET_0_73460);
    
    HIEFFPLA_INST_0_55464 : OA1C
      port map(A => HIEFFPLA_NET_0_75511, B => 
        HIEFFPLA_NET_0_75510, C => 
        \Communications_0/UART_0/tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75505);
    
    HIEFFPLA_INST_0_70335 : AOI1D
      port map(A => General_Controller_0_st_ren1, B => 
        \SweepTable_0/WEBP\, C => 
        \General_Controller_0_st_raddr_1[0]\, Y => 
        \TableSelect_0_RADDR[0]\);
    
    HIEFFPLA_INST_0_69961 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        B => HIEFFPLA_NET_0_72228, C => HIEFFPLA_NET_0_72231, Y
         => HIEFFPLA_NET_0_72259);
    
    \Science_0/ADC_READ_0/cnt1dn[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73402, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1dn[6]_net_1\);
    
    HIEFFPLA_INST_0_67652 : AOI1
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72833);
    
    HIEFFPLA_INST_0_68388 : AOI1
      port map(A => HIEFFPLA_NET_0_72671, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[7]\, C => 
        HIEFFPLA_NET_0_72659, Y => HIEFFPLA_NET_0_72660);
    
    HIEFFPLA_INST_0_70464 : AND3
      port map(A => \Timekeeper_0_milliseconds[15]\, B => 
        HIEFFPLA_NET_0_72118, C => 
        \Timekeeper_0_milliseconds[16]\, Y => 
        HIEFFPLA_NET_0_72121);
    
    HIEFFPLA_INST_0_61123 : NOR3A
      port map(A => \General_Controller_0/command[1]_net_1\, B
         => \General_Controller_0/command[4]_net_1\, C => 
        \General_Controller_0/command[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74271);
    
    HIEFFPLA_INST_0_69652 : AO1
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        B => PRESSURE_SCL_c, C => HIEFFPLA_NET_0_72341, Y => 
        HIEFFPLA_NET_0_72336);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRY[2]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75314, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[2]\\\\\);
    
    HIEFFPLA_INST_0_58338 : AO1
      port map(A => \Sensors_0_acc_x[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74797, Y => HIEFFPLA_NET_0_74798);
    
    \Timing_0/m_time[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72061, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_time[4]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[68]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[12]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[68]\);
    
    HIEFFPLA_INST_0_66969 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[0]\, 
        B => \Sensors_0/Accelerometer_0/state[8]\, C => 
        HIEFFPLA_NET_0_72986, Y => HIEFFPLA_NET_0_72995);
    
    HIEFFPLA_INST_0_69061 : AND2B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72481);
    
    HIEFFPLA_INST_0_67259 : AND3
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72925);
    
    \FMC_DA_pad[2]/U0/U1\ : IOTRI_OB_EB
      port map(D => \FMC_DA_c[2]\, E => \VCC\, DOUT => 
        \FMC_DA_pad[2]/U0/NET1\, EOUT => \FMC_DA_pad[2]/U0/NET2\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[10]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72782, Q => 
        \Sensors_0_mag_y[10]\);
    
    HIEFFPLA_INST_0_64711 : AO1A
      port map(A => 
        \General_Controller_0/uc_tx_substate[2]_net_1\, B => 
        HIEFFPLA_NET_0_73553, C => HIEFFPLA_NET_0_73554, Y => 
        HIEFFPLA_NET_0_73555);
    
    HIEFFPLA_INST_0_67477 : AO1A
      port map(A => HIEFFPLA_NET_0_72836, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_72943, Y => HIEFFPLA_NET_0_72869);
    
    HIEFFPLA_INST_0_63800 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[4]_net_1\, 
        B => \General_Controller_0/sweep_table_points[4]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73709);
    
    HIEFFPLA_INST_0_60134 : AO1A
      port map(A => HIEFFPLA_NET_0_74638, B => 
        \GS_Readout_0/subState[1]_net_1\, C => 
        HIEFFPLA_NET_0_74616, Y => HIEFFPLA_NET_0_74456);
    
    HIEFFPLA_INST_0_68749 : AO1A
      port map(A => GYRO_SCL_c, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, C => 
        HIEFFPLA_NET_0_72629, Y => HIEFFPLA_NET_0_72571);
    
    HIEFFPLA_INST_0_61816 : XA1B
      port map(A => 
        \General_Controller_0/sweep_table_write_wait[0]_net_1\, B
         => HIEFFPLA_NET_0_74127, C => HIEFFPLA_NET_0_73806, Y
         => HIEFFPLA_NET_0_74123);
    
    \General_Controller_0/uc_rx_state[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73867, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_state[4]_net_1\);
    
    HIEFFPLA_INST_0_71119 : AOI1D
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => \Sensors_0_acc_temp[0]\, Y => HIEFFPLA_NET_0_71979);
    
    HIEFFPLA_INST_0_70638 : XA1B
      port map(A => \Timing_0/s_count[0]_net_1\, B => 
        HIEFFPLA_NET_0_72083, C => HIEFFPLA_NET_0_72058, Y => 
        HIEFFPLA_NET_0_72056);
    
    HIEFFPLA_INST_0_71084 : AO1A
      port map(A => Communications_0_ext_tx_rdy, B => 
        HIEFFPLA_NET_0_71981, C => HIEFFPLA_NET_0_74610, Y => 
        HIEFFPLA_NET_0_74611);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[21]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[21]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[21]\);
    
    HIEFFPLA_INST_0_56036 : XA1A
      port map(A => HIEFFPLA_NET_0_75276, B => 
        HIEFFPLA_NET_0_75331, C => HIEFFPLA_NET_0_75362, Y => 
        HIEFFPLA_NET_0_75363);
    
    HIEFFPLA_INST_0_55350 : AND2B
      port map(A => HIEFFPLA_NET_0_75529, B => 
        \Communications_0/UART_0/tx_clk_count_i_0[5]\, Y => 
        HIEFFPLA_NET_0_75534);
    
    HIEFFPLA_INST_0_70097 : NOR3B
      port map(A => HIEFFPLA_NET_0_72209, B => 
        HIEFFPLA_NET_0_72286, C => HIEFFPLA_NET_0_72273, Y => 
        HIEFFPLA_NET_0_72219);
    
    HIEFFPLA_INST_0_60922 : NOR2A
      port map(A => HIEFFPLA_NET_0_74318, B => 
        \General_Controller_0/un10_uc_tx_rdy_i[4]\, Y => 
        HIEFFPLA_NET_0_74319);
    
    HIEFFPLA_INST_0_70166 : NAND3B
      port map(A => HIEFFPLA_NET_0_72197, B => 
        HIEFFPLA_NET_0_72179, C => HIEFFPLA_NET_0_72203, Y => 
        HIEFFPLA_NET_0_72204);
    
    HIEFFPLA_INST_0_58648 : NAND3C
      port map(A => HIEFFPLA_NET_0_74701, B => 
        HIEFFPLA_NET_0_74646, C => HIEFFPLA_NET_0_74621, Y => 
        HIEFFPLA_NET_0_74713);
    
    HIEFFPLA_INST_0_57146 : AND2
      port map(A => \ch3_data_net_0[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75154);
    
    HIEFFPLA_INST_0_66730 : NAND2B
      port map(A => ACCE_SCL_c, B => HIEFFPLA_NET_0_73144, Y => 
        HIEFFPLA_NET_0_73052);
    
    HIEFFPLA_INST_0_61581 : AND3
      port map(A => HIEFFPLA_NET_0_73777, B => 
        HIEFFPLA_NET_0_74172, C => HIEFFPLA_NET_0_73918, Y => 
        HIEFFPLA_NET_0_74179);
    
    HIEFFPLA_INST_0_58409 : AND2
      port map(A => HIEFFPLA_NET_0_74771, B => 
        \Data_Saving_0/Packet_Saver_0/gyro_flag_net_1\, Y => 
        HIEFFPLA_NET_0_74775);
    
    \General_Controller_0/sweep_table_step_id[7]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73926, Q => 
        \General_Controller_0/sweep_table_step_id[7]_net_1\);
    
    \Timing_0/s_time[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72044, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_time[1]_net_1\);
    
    HIEFFPLA_INST_0_69403 : NOR3B
      port map(A => HIEFFPLA_NET_0_72351, B => 
        HIEFFPLA_NET_0_72373, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72397);
    
    HIEFFPLA_INST_0_55839 : NAND3C
      port map(A => \Communications_0/UART_1/tx_clk_count_i_0[6]\, 
        B => \Communications_0/UART_1/tx_clk_count_i_0[5]\, C => 
        HIEFFPLA_NET_0_75412, Y => HIEFFPLA_NET_0_75414);
    
    HIEFFPLA_INST_0_64145 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_1[3]_net_1\, 
        B => 
        \General_Controller_0/constant_bias_voltage_1[11]_net_1\, 
        S => \General_Controller_0/uc_tx_substate[1]_net_1\, Y
         => HIEFFPLA_NET_0_73662);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72216, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\);
    
    HIEFFPLA_INST_0_58460 : MX2C
      port map(A => HIEFFPLA_NET_0_74759, B => 
        HIEFFPLA_NET_0_74754, S => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74761);
    
    HIEFFPLA_INST_0_61132 : AO1
      port map(A => Pressure_Signal_Debounce_0_low_pressure, B
         => \General_Controller_0/flight_state[3]_net_1\, C => 
        \General_Controller_0/mission_mode_net_1\, Y => 
        HIEFFPLA_NET_0_74269);
    
    \Science_0/ADC_READ_0/g2i[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73259, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73420, Q => 
        \Science_0/ADC_READ_0_G2[1]\);
    
    HIEFFPLA_INST_0_60835 : NOR2A
      port map(A => HIEFFPLA_NET_0_74636, B => 
        HIEFFPLA_NET_0_74382, Y => HIEFFPLA_NET_0_74349);
    
    HIEFFPLA_INST_0_60116 : NOR2A
      port map(A => HIEFFPLA_NET_0_74380, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74459);
    
    \Science_0/ADC_READ_0/exp_packet_1[60]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[4]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[60]\);
    
    \RESET_pad/U0/U1\ : IOIN_IB
      port map(YIN => \RESET_pad/U0/NET1\, Y => RESET_c);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[9]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72281, Q => \Sensors_0_pressure_raw[9]\);
    
    HIEFFPLA_INST_0_66190 : AO1
      port map(A => \Science_0/SET_LP_GAIN_0/state[5]_net_1\, B
         => \Science_0/ADC_READ_0_G3[0]\, C => 
        HIEFFPLA_NET_0_73163, Y => HIEFFPLA_NET_0_73183);
    
    HIEFFPLA_INST_0_58967 : NOR3B
      port map(A => Communications_0_ext_tx_rdy, B => 
        \GS_Readout_0/state[5]_net_1\, C => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74647);
    
    \General_Controller_0/ext_oen\ : DFN1E1C1
      port map(D => Communications_0_ext_rx_rdy, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74302, Q => General_Controller_0_ext_oen);
    
    \Science_0/ADC_READ_0/data_a[8]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[8]_net_1\);
    
    HIEFFPLA_INST_0_64445 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state_0[4]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[0]_net_1\, C => 
        HIEFFPLA_NET_0_73875, Y => HIEFFPLA_NET_0_73625);
    
    HIEFFPLA_INST_0_57204 : AO1
      port map(A => \Sensors_0_pressure_time[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75090, Y => HIEFFPLA_NET_0_75131);
    
    HIEFFPLA_INST_0_70783 : AOI1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72013);
    
    HIEFFPLA_INST_0_68074 : OR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72739);
    
    HIEFFPLA_INST_0_64247 : MX2
      port map(A => HIEFFPLA_NET_0_73741, B => 
        HIEFFPLA_NET_0_73733, S => HIEFFPLA_NET_0_73588, Y => 
        HIEFFPLA_NET_0_73645);
    
    HIEFFPLA_INST_0_66352 : OR3A
      port map(A => HIEFFPLA_NET_0_73139, B => 
        HIEFFPLA_NET_0_73060, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_73140);
    
    \General_Controller_0/sweep_table_samples_per_step[8]\ : 
        DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[0]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[8]_net_1\);
    
    \Communications_0/UART_1/tx_clk_count[5]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75406, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_clk_count_i_0[5]\);
    
    HIEFFPLA_INST_0_69046 : NOR3A
      port map(A => HIEFFPLA_NET_0_72478, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72486);
    
    HIEFFPLA_INST_0_63284 : OR2A
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_substate[2]_net_1\, Y
         => HIEFFPLA_NET_0_73788);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/state[8]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73061, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/state[8]\);
    
    HIEFFPLA_INST_0_66473 : OA1C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\, 
        B => HIEFFPLA_NET_0_73113, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_73111);
    
    \Timing_0/f_time[0]\ : DFN1C1
      port map(D => \AFLSDF_INV_9\, CLK => CLKINT_0_Y_0, CLR => 
        CLKINT_1_Y, Q => \Timing_0/f_time[0]_net_1\);
    
    HIEFFPLA_INST_0_61879 : NOR3A
      port map(A => \General_Controller_0/uc_rx_byte[4]_net_1\, B
         => HIEFFPLA_NET_0_74109, C => HIEFFPLA_NET_0_74084, Y
         => HIEFFPLA_NET_0_74110);
    
    HIEFFPLA_INST_0_56325 : XOR2
      port map(A => HIEFFPLA_NET_0_75294, B => 
        HIEFFPLA_NET_0_75312, Y => HIEFFPLA_NET_0_75310);
    
    HIEFFPLA_INST_0_62542 : NAND3C
      port map(A => HIEFFPLA_NET_0_73797, B => 
        HIEFFPLA_NET_0_74023, C => HIEFFPLA_NET_0_73866, Y => 
        HIEFFPLA_NET_0_73960);
    
    HIEFFPLA_INST_0_64621 : AND3B
      port map(A => HIEFFPLA_NET_0_73977, B => 
        HIEFFPLA_NET_0_73928, C => HIEFFPLA_NET_0_73583, Y => 
        HIEFFPLA_NET_0_73584);
    
    HIEFFPLA_INST_0_58795 : AND2
      port map(A => \General_Controller_0_gs_id[3]\, B => 
        HIEFFPLA_NET_0_74484, Y => HIEFFPLA_NET_0_74683);
    
    HIEFFPLA_INST_0_63770 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[7]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[7]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73714);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73067, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_net_1\);
    
    HIEFFPLA_INST_0_68636 : AND2
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, B => 
        GYRO_SCL_c, Y => HIEFFPLA_NET_0_72600);
    
    \Science_0/ADC_READ_0/chan6_data[0]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[0]\);
    
    \Science_0/ADC_READ_0/chan0_data[0]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[0]\);
    
    HIEFFPLA_INST_0_68233 : NOR3B
      port map(A => HIEFFPLA_NET_0_72702, B => 
        HIEFFPLA_NET_0_72626, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_72699);
    
    HIEFFPLA_INST_0_56008 : NAND3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[2]\\\\\, B
         => HIEFFPLA_NET_0_75308, C => 
        \Data_Saving_0/Packet_Saver_0_we\, Y => 
        HIEFFPLA_NET_0_75370);
    
    HIEFFPLA_INST_0_61955 : AO1
      port map(A => HIEFFPLA_NET_0_73791, B => 
        HIEFFPLA_NET_0_74026, C => HIEFFPLA_NET_0_74089, Y => 
        HIEFFPLA_NET_0_74090);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRY[10]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75267, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[10]\\\\\);
    
    HIEFFPLA_INST_0_70495 : XOR2
      port map(A => HIEFFPLA_NET_0_72118, B => 
        \Timekeeper_0_milliseconds[15]\, Y => 
        HIEFFPLA_NET_0_72110);
    
    HIEFFPLA_INST_0_57133 : AO1
      port map(A => \Sensors_0_pressure_time[14]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75101, Y => HIEFFPLA_NET_0_75163);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[10]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72490, Q => 
        \ch3_data_net_0[6]\);
    
    HIEFFPLA_INST_0_65680 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt4dn[7]_net_1\, B => 
        HIEFFPLA_NET_0_73310, C => HIEFFPLA_NET_0_73274, Y => 
        HIEFFPLA_NET_0_73311);
    
    \General_Controller_0/unit_id[7]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73990, Q => 
        \General_Controller_0_unit_id[7]\);
    
    HIEFFPLA_INST_0_55827 : AOI1C
      port map(A => \Communications_0/UART_1/tx_state[0]_net_1\, 
        B => \Communications_0/UART_1/tx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_75420, Y => HIEFFPLA_NET_0_75419);
    
    HIEFFPLA_INST_0_55848 : NAND3C
      port map(A => HIEFFPLA_NET_0_75418, B => 
        \Communications_0/UART_1/tx_clk_count_i_0[3]\, C => 
        \Communications_0/UART_1/tx_clk_count_i_0[4]\, Y => 
        HIEFFPLA_NET_0_75412);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[2]\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72406, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72352, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[2]_net_1\);
    
    HIEFFPLA_INST_0_66290 : AO1C
      port map(A => HIEFFPLA_NET_0_73175, B => 
        \Science_0/SET_LP_GAIN_0/state[6]_net_1\, C => 
        \Science_0/SET_LP_GAIN_0/state_i_0[2]\, Y => 
        HIEFFPLA_NET_0_73154);
    
    HIEFFPLA_INST_0_56347 : AX1C
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[6]\\\\\, B
         => HIEFFPLA_NET_0_75348, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[7]\\\\\, Y
         => HIEFFPLA_NET_0_75304);
    
    HIEFFPLA_INST_0_56400 : XOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, B
         => HIEFFPLA_NET_0_75352, C => HIEFFPLA_NET_0_75262, Y
         => HIEFFPLA_NET_0_75289);
    
    HIEFFPLA_INST_0_61911 : AND3C
      port map(A => HIEFFPLA_NET_0_74100, B => 
        \General_Controller_0/uc_rx_byte[0]_net_1\, C => 
        \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74101);
    
    AFLSDF_INV_21 : INV
      port map(A => \ClockDivs_0/cnt_800kHz[0]_net_1\, Y => 
        \AFLSDF_INV_21\);
    
    \Science_0/ADC_READ_0/chan5_data[8]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[8]\);
    
    \General_Controller_0/sweep_table_read_wait[30]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74152, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/sweep_table_read_wait[30]_net_1\);
    
    HIEFFPLA_INST_0_56364 : AX1D
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, B
         => HIEFFPLA_NET_0_75371, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\, Y
         => HIEFFPLA_NET_0_75300);
    
    \Science_0/ADC_READ_0/chan2_data[11]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[17]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[11]\);
    
    HIEFFPLA_INST_0_68719 : AOI1
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\, B
         => \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_72579);
    
    HIEFFPLA_INST_0_66130 : NOR2A
      port map(A => \Science_0/DAC_SET_0/vector[13]_net_1\, B => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73199);
    
    HIEFFPLA_INST_0_70344 : AOI1D
      port map(A => General_Controller_0_st_ren1, B => 
        \SweepTable_0/WEBP\, C => 
        \General_Controller_0_st_raddr_1[4]\, Y => 
        \TableSelect_0_RADDR[4]\);
    
    \Science_0/ADC_READ_0/g4i[0]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73250, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73421, Q => 
        \Science_0/ADC_READ_0_G4[0]\);
    
    HIEFFPLA_INST_0_66576 : MX2
      port map(A => HIEFFPLA_NET_0_73087, B => 
        HIEFFPLA_NET_0_73086, S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73089);
    
    HIEFFPLA_INST_0_66728 : AND2B
      port map(A => HIEFFPLA_NET_0_73142, B => 
        \Sensors_0/Accelerometer_0/state[8]\, Y => 
        HIEFFPLA_NET_0_73053);
    
    \General_Controller_0/sweep_table_samples_per_step[1]\ : 
        DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[1]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[1]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRYSYNC[4]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_4_Q\, CLK
         => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[4]\\\\\);
    
    \General_Controller_0/uc_rx_state_0[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73895, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\);
    
    HIEFFPLA_INST_0_57471 : AO1
      port map(A => \Sensors_0_acc_z[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74863, Y => HIEFFPLA_NET_0_75036);
    
    HIEFFPLA_INST_0_69684 : OR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[2]_net_1\, 
        B => HIEFFPLA_NET_0_72381, C => HIEFFPLA_NET_0_72388, Y
         => HIEFFPLA_NET_0_72330);
    
    HIEFFPLA_INST_0_61011 : NAND2
      port map(A => \General_Controller_0/flight_state[3]_net_1\, 
        B => \General_Controller_0/mission_mode_net_1\, Y => 
        HIEFFPLA_NET_0_74296);
    
    HIEFFPLA_INST_0_68012 : NOR3B
      port map(A => HIEFFPLA_NET_0_72738, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        C => HIEFFPLA_NET_0_72939, Y => HIEFFPLA_NET_0_72754);
    
    \Science_0/ADC_READ_0/cnt4dn[5]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73313, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4dn[5]_net_1\);
    
    HIEFFPLA_INST_0_56227 : XOR2
      port map(A => HIEFFPLA_NET_0_75323, B => 
        HIEFFPLA_NET_0_75322, Y => HIEFFPLA_NET_0_75330);
    
    HIEFFPLA_INST_0_65263 : AND3B
      port map(A => \Sensors_0_pressure_raw[5]\, B => 
        \Sensors_0_pressure_raw[1]\, C => HIEFFPLA_NET_0_73469, Y
         => HIEFFPLA_NET_0_73431);
    
    HIEFFPLA_INST_0_57433 : AO1
      port map(A => \Sensors_0_acc_z[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74868, Y => HIEFFPLA_NET_0_75047);
    
    HIEFFPLA_INST_0_67782 : AND3C
      port map(A => HIEFFPLA_NET_0_72765, B => 
        HIEFFPLA_NET_0_72903, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72803);
    
    \Science_0/ADC_READ_0/cnt4dn[4]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73314, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4dn[4]_net_1\);
    
    \General_Controller_0/sweep_table_read_value[14]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74165, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[14]_net_1\);
    
    \Timekeeper_0/milliseconds[12]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72113, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[12]\);
    
    HIEFFPLA_INST_0_63930 : AND2
      port map(A => HIEFFPLA_NET_0_73659, B => 
        HIEFFPLA_NET_0_73594, Y => HIEFFPLA_NET_0_73688);
    
    HIEFFPLA_INST_0_69864 : AO1B
      port map(A => HIEFFPLA_NET_0_72223, B => 
        Sensors_0_pressure_new_data, C => HIEFFPLA_NET_0_72241, Y
         => HIEFFPLA_NET_0_72287);
    
    \General_Controller_0/sweep_table_sweep_cnt[12]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74141, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[12]_net_1\);
    
    \GS_Readout_0/subState[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74351, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/subState[4]_net_1\);
    
    \TOP_UART_TX_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => SCIENCE_TX_c_c, E => \VCC\, DOUT => 
        \TOP_UART_TX_pad/U0/NET1\, EOUT => 
        \TOP_UART_TX_pad/U0/NET2\);
    
    \LED1_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => LED1_c, E => \VCC\, DOUT => 
        \LED1_pad/U0/NET1\, EOUT => \LED1_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_58054 : AO1
      port map(A => \Sensors_0_gyro_y[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75161, Y => HIEFFPLA_NET_0_74868);
    
    HIEFFPLA_INST_0_69736 : AX1
      port map(A => HIEFFPLA_NET_0_72394, B => 
        HIEFFPLA_NET_0_72380, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72319);
    
    HIEFFPLA_INST_0_57284 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[42]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75096);
    
    HIEFFPLA_INST_0_69326 : XO1
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => HIEFFPLA_NET_0_72321, C => HIEFFPLA_NET_0_72415, Y
         => HIEFFPLA_NET_0_72418);
    
    HIEFFPLA_INST_0_64866 : NAND3C
      port map(A => HIEFFPLA_NET_0_73616, B => 
        HIEFFPLA_NET_0_73555, C => HIEFFPLA_NET_0_73613, Y => 
        HIEFFPLA_NET_0_73522);
    
    HIEFFPLA_INST_0_62101 : AO1A
      port map(A => HIEFFPLA_NET_0_73890, B => 
        HIEFFPLA_NET_0_73906, C => HIEFFPLA_NET_0_74051, Y => 
        HIEFFPLA_NET_0_74052);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[2]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_75251, CLK => CLKINT_0_Y_0, E
         => CLKINT_1_Y, Q => 
        \Data_Saving_0/Interrupt_Generator_0/counter[2]_net_1\);
    
    HIEFFPLA_INST_0_61008 : NAND2B
      port map(A => \General_Controller_0/flight_state[0]_net_1\, 
        B => \General_Controller_0/flight_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74297);
    
    HIEFFPLA_INST_0_59265 : MX2
      port map(A => HIEFFPLA_NET_0_74442, B => 
        HIEFFPLA_NET_0_74431, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74577);
    
    HIEFFPLA_INST_0_70530 : XOR2
      port map(A => HIEFFPLA_NET_0_72124, B => 
        \Timekeeper_0_milliseconds[9]\, Y => HIEFFPLA_NET_0_72093);
    
    HIEFFPLA_INST_0_70975 : AO1B
      port map(A => \Science_0/ADC_READ_0/cnt4up[4]_net_1\, B => 
        HIEFFPLA_NET_0_73276, C => \Science_0/ADC_READ_0_G4[0]\, 
        Y => HIEFFPLA_NET_0_71996);
    
    \Science_0/ADC_READ_0/exp_new_data\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/newflag_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73273, Q => Science_0_exp_new_data);
    
    HIEFFPLA_INST_0_70777 : XA1A
      port map(A => HIEFFPLA_NET_0_72014, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[7]_net_1\, 
        C => HIEFFPLA_NET_0_72236, Y => HIEFFPLA_NET_0_72292);
    
    HIEFFPLA_INST_0_58988 : OR3A
      port map(A => HIEFFPLA_NET_0_74638, B => 
        \GS_Readout_0/state[0]_net_1\, C => 
        \GS_Readout_0/state[6]_net_1\, Y => HIEFFPLA_NET_0_74643);
    
    \General_Controller_0/constant_bias_voltage_0[1]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[1]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[1]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[7]\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72292, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72221, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[7]_net_1\);
    
    HIEFFPLA_INST_0_67637 : OR2A
      port map(A => HIEFFPLA_NET_0_72798, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, Y
         => HIEFFPLA_NET_0_72836);
    
    HIEFFPLA_INST_0_63170 : NAND3C
      port map(A => HIEFFPLA_NET_0_73796, B => 
        HIEFFPLA_NET_0_73804, C => HIEFFPLA_NET_0_73958, Y => 
        HIEFFPLA_NET_0_73816);
    
    HIEFFPLA_INST_0_64962 : AX1C
      port map(A => HIEFFPLA_NET_0_73501, B => 
        \I2C_PassThrough_0/cnt[2]_net_1\, C => 
        \I2C_PassThrough_0/cnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73502);
    
    \Science_0/ADC_READ_0/exp_packet_1[1]\ : DFN1E0
      port map(D => \AFLSDF_INV_10\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[1]\);
    
    HIEFFPLA_INST_0_70764 : OA1C
      port map(A => HIEFFPLA_NET_0_72017, B => 
        HIEFFPLA_NET_0_72286, C => HIEFFPLA_NET_0_72018, Y => 
        HIEFFPLA_NET_0_72178);
    
    HIEFFPLA_INST_0_67635 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72837);
    
    HIEFFPLA_INST_0_62117 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state_0[1]_net_1\, 
        B => HIEFFPLA_NET_0_73888, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74049);
    
    HIEFFPLA_INST_0_64593 : AND2B
      port map(A => \General_Controller_0/uc_tx_state[3]_net_1\, 
        B => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73593);
    
    \General_Controller_0/uc_rx_substate[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73770, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_substate[4]_net_1\);
    
    \Timing_0/m_time[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72064, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_time[1]_net_1\);
    
    HIEFFPLA_INST_0_65004 : XA1
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[4]_net_1\, 
        B => HIEFFPLA_NET_0_73444, C => HIEFFPLA_NET_0_73490, Y
         => HIEFFPLA_NET_0_73491);
    
    HIEFFPLA_INST_0_60603 : XA1
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, C => 
        HIEFFPLA_NET_0_74365, Y => HIEFFPLA_NET_0_74389);
    
    \General_Controller_0/uc_rx_byte[6]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[6]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte[6]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[7]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72753, Q => 
        \Sensors_0_acc_z[7]\);
    
    \General_Controller_0/constant_bias_probe_id[4]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73923, Q => 
        \General_Controller_0/un10_uc_tx_rdy_i[4]\);
    
    HIEFFPLA_INST_0_67178 : AND3
      port map(A => HIEFFPLA_NET_0_72957, B => 
        HIEFFPLA_NET_0_72954, C => HIEFFPLA_NET_0_72951, Y => 
        HIEFFPLA_NET_0_72945);
    
    HIEFFPLA_INST_0_67457 : XO1A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        C => HIEFFPLA_NET_0_72873, Y => HIEFFPLA_NET_0_72874);
    
    HIEFFPLA_INST_0_64427 : MX2
      port map(A => HIEFFPLA_NET_0_73707, B => 
        HIEFFPLA_NET_0_73699, S => HIEFFPLA_NET_0_73593, Y => 
        HIEFFPLA_NET_0_73627);
    
    HIEFFPLA_INST_0_69983 : NOR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_s_ack_error\, Y
         => HIEFFPLA_NET_0_72253);
    
    \Timekeeper_0/milliseconds[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72105, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[1]\);
    
    \General_Controller_0/sweep_table_sample_skip[2]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[2]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[2]_net_1\);
    
    HIEFFPLA_INST_0_55817 : MX2C
      port map(A => \Communications_0/UART_1/tx_byte[3]_net_1\, B
         => \Communications_0/UART_1/tx_byte[7]_net_1\, S => 
        \Communications_0/UART_1/tx_count[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75421);
    
    HIEFFPLA_INST_0_62818 : NOR3A
      port map(A => HIEFFPLA_NET_0_74014, B => 
        HIEFFPLA_NET_0_73813, C => HIEFFPLA_NET_0_73899, Y => 
        HIEFFPLA_NET_0_73894);
    
    HIEFFPLA_INST_0_62518 : AND3
      port map(A => HIEFFPLA_NET_0_74029, B => 
        HIEFFPLA_NET_0_73921, C => HIEFFPLA_NET_0_73780, Y => 
        HIEFFPLA_NET_0_73966);
    
    HIEFFPLA_INST_0_55039 : NOR3B
      port map(A => HIEFFPLA_NET_0_75599, B => 
        HIEFFPLA_NET_0_75604, C => 
        \Communications_0/UART_0/rx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75607);
    
    HIEFFPLA_INST_0_64189 : NOR3A
      port map(A => HIEFFPLA_NET_0_73749, B => 
        \General_Controller_0/uc_tx_state[12]_net_1\, C => 
        \General_Controller_0/uc_tx_state[14]_net_1\, Y => 
        HIEFFPLA_NET_0_73653);
    
    \General_Controller_0/constant_bias_probe_id[6]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73923, Q => 
        \General_Controller_0/un10_uc_tx_rdy_i[6]\);
    
    HIEFFPLA_INST_0_65038 : XOR2
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[0]_net_1\, 
        B => HIEFFPLA_NET_0_73478, Y => HIEFFPLA_NET_0_73483);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1E1C0_data_out[1]\\\\/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75286, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \FMC_DA_c[1]\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRYSYNC[5]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_18_Q\, 
        CLK => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[5]\\\\\);
    
    HIEFFPLA_INST_0_62702 : AND3
      port map(A => HIEFFPLA_NET_0_73883, B => 
        HIEFFPLA_NET_0_73887, C => HIEFFPLA_NET_0_73775, Y => 
        HIEFFPLA_NET_0_73925);
    
    HIEFFPLA_INST_0_66879 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_we\, 
        B => \Sensors_0/Accelerometer_0/state[8]\, Y => 
        HIEFFPLA_NET_0_73013);
    
    HIEFFPLA_INST_0_59119 : AO1A
      port map(A => HIEFFPLA_NET_0_74592, B => 
        \GS_Readout_0/prevState[2]_net_1\, C => 
        HIEFFPLA_NET_0_74586, Y => HIEFFPLA_NET_0_74608);
    
    \General_Controller_0/gs_id[0]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73922, Q => 
        \General_Controller_0_gs_id[0]\);
    
    HIEFFPLA_INST_0_65296 : NOR3B
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, B => 
        \Science_0/ADC_READ_0/newflag_net_1\, C => 
        \Science_0/ADC_READ_0/chan[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73419);
    
    \Eject_Signal_Debounce_0/ms_cnt[4]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74742, CLK => CLKINT_0_Y_0, Q
         => \Eject_Signal_Debounce_0/ms_cnt[4]_net_1\);
    
    HIEFFPLA_INST_0_68335 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, B => 
        HIEFFPLA_NET_0_72678, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_72679);
    
    HIEFFPLA_INST_0_67517 : NAND3C
      port map(A => HIEFFPLA_NET_0_72858, B => 
        HIEFFPLA_NET_0_72849, C => HIEFFPLA_NET_0_72818, Y => 
        HIEFFPLA_NET_0_72859);
    
    HIEFFPLA_INST_0_67440 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, Y
         => HIEFFPLA_NET_0_72879);
    
    HIEFFPLA_INST_0_70369 : AND3
      port map(A => \Timekeeper_0_microseconds[17]\, B => 
        HIEFFPLA_NET_0_72162, C => 
        \Timekeeper_0_microseconds[18]\, Y => 
        HIEFFPLA_NET_0_72158);
    
    HIEFFPLA_INST_0_56005 : NOR2A
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, B
         => HIEFFPLA_NET_0_75370, Y => HIEFFPLA_NET_0_75371);
    
    \Science_0/ADC_READ_0/chan7_data[0]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[0]\);
    
    HIEFFPLA_INST_0_65327 : AND2B
      port map(A => \Science_0/ADC_READ_0/cnt1dn[0]_net_1\, B => 
        HIEFFPLA_NET_0_73244, Y => HIEFFPLA_NET_0_73408);
    
    HIEFFPLA_INST_0_60853 : AX1B
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, C => 
        \GS_Readout_0/subState[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74341);
    
    HIEFFPLA_INST_0_58712 : NOR3B
      port map(A => HIEFFPLA_NET_0_74641, B => 
        HIEFFPLA_NET_0_74499, C => HIEFFPLA_NET_0_74552, Y => 
        HIEFFPLA_NET_0_74699);
    
    HIEFFPLA_INST_0_58374 : AND2
      port map(A => \Sensors_0_mag_z[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        Y => HIEFFPLA_NET_0_74788);
    
    HIEFFPLA_INST_0_70955 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[0]\, 
        C => HIEFFPLA_NET_0_72884, Y => HIEFFPLA_NET_0_72002);
    
    \Timing_0/m_count[7]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72028, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_count[7]_net_1\);
    
    HIEFFPLA_INST_0_67542 : AO1
      port map(A => HIEFFPLA_NET_0_72848, B => 
        HIEFFPLA_NET_0_72830, C => HIEFFPLA_NET_0_72822, Y => 
        HIEFFPLA_NET_0_72856);
    
    HIEFFPLA_INST_0_57765 : AO1B
      port map(A => \Data_Hub_Packets_0_status_packet[63]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, C
         => HIEFFPLA_NET_0_74948, Y => HIEFFPLA_NET_0_74949);
    
    HIEFFPLA_INST_0_58266 : AO1
      port map(A => \Sensors_0_gyro_x[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74815, Y => HIEFFPLA_NET_0_74816);
    
    \GYRO_SCL_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => GYRO_SCL_c, E => \VCC\, DOUT => 
        \GYRO_SCL_pad/U0/NET1\, EOUT => \GYRO_SCL_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_62181 : AO1E
      port map(A => HIEFFPLA_NET_0_73915, B => 
        HIEFFPLA_NET_0_73973, C => HIEFFPLA_NET_0_73775, Y => 
        HIEFFPLA_NET_0_74035);
    
    HIEFFPLA_INST_0_55635 : XA1A
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[28]_net_1\, B => 
        HIEFFPLA_NET_0_75467, C => HIEFFPLA_NET_0_75437, Y => 
        HIEFFPLA_NET_0_75459);
    
    HIEFFPLA_INST_0_55873 : NAND2B
      port map(A => HIEFFPLA_NET_0_75399, B => 
        HIEFFPLA_NET_0_75419, Y => HIEFFPLA_NET_0_75407);
    
    HIEFFPLA_INST_0_63602 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[11]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_sample_skip[11]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73742);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[22]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[22]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[22]\);
    
    HIEFFPLA_INST_0_63542 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[9]_net_1\, B
         => \General_Controller_0/sweep_table_points[9]_net_1\, S
         => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73752);
    
    \Science_0/ADC_READ_0/cnt3up[0]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73336, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3up[0]_net_1\);
    
    HIEFFPLA_INST_0_71218 : MIN3X
      port map(A => 
        \Communications_0/FFU_Command_Checker_0/state[0]_net_1\, 
        B => 
        \Communications_0/FFU_Command_Checker_0/state[1]_net_1\, 
        C => \Communications_0/UART_0_rx_rdy\, Y => 
        HIEFFPLA_NET_0_71970);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_72469, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\);
    
    HIEFFPLA_INST_0_56118 : XNOR3
      port map(A => HIEFFPLA_NET_0_75321, B => 
        HIEFFPLA_NET_0_75288, C => HIEFFPLA_NET_0_75324, Y => 
        HIEFFPLA_NET_0_75343);
    
    \Communications_0/UART_0/tx\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75544, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => \Communications_0/UART_0_tx\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[1]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[1]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[1]\);
    
    HIEFFPLA_INST_0_65365 : AND2
      port map(A => \Science_0/ADC_READ_0/cnt1dn[5]_net_1\, B => 
        HIEFFPLA_NET_0_73413, Y => HIEFFPLA_NET_0_73398);
    
    HIEFFPLA_INST_0_57529 : AO1B
      port map(A => \Sensors_0_mag_z[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75018, Y => HIEFFPLA_NET_0_75019);
    
    HIEFFPLA_INST_0_70266 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        B => \Sensors_0/Pressure_Sensor_0/state[8]\, C => 
        HIEFFPLA_NET_0_72269, Y => HIEFFPLA_NET_0_72183);
    
    HIEFFPLA_INST_0_63794 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[3]_net_1\, 
        B => \General_Controller_0/sweep_table_points[3]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73710);
    
    HIEFFPLA_INST_0_63209 : NOR3B
      port map(A => HIEFFPLA_NET_0_73918, B => 
        \General_Controller_0/uc_rx_substate[3]_net_1\, C => 
        HIEFFPLA_NET_0_73782, Y => HIEFFPLA_NET_0_73806);
    
    HIEFFPLA_INST_0_60824 : XA1B
      port map(A => HIEFFPLA_NET_0_74346, B => 
        \GS_Readout_0/subState[3]_net_1\, C => 
        HIEFFPLA_NET_0_74350, Y => HIEFFPLA_NET_0_74352);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/data_out_1[0]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_72570, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72547, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[0]\);
    
    HIEFFPLA_INST_0_68422 : MX2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[2]\, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[6]\, S => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72654);
    
    HIEFFPLA_INST_0_64061 : MX2
      port map(A => HIEFFPLA_NET_0_73638, B => 
        HIEFFPLA_NET_0_73630, S => HIEFFPLA_NET_0_73585, Y => 
        HIEFFPLA_NET_0_73675);
    
    \Science_0/ADC_READ_0/exp_packet_1[62]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[6]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[62]\);
    
    HIEFFPLA_INST_0_67514 : AND2
      port map(A => HIEFFPLA_NET_0_72778, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72860);
    
    \General_Controller_0/sweep_table_points[12]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[12]_net_1\);
    
    AFLSDF_INV_37 : INV
      port map(A => CLKINT_1_Y, Y => \AFLSDF_INV_37\);
    
    HIEFFPLA_INST_0_65542 : NOR2A
      port map(A => HIEFFPLA_NET_0_73349, B => 
        \Science_0/ADC_READ_0/cnt3dn[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73347);
    
    HIEFFPLA_INST_0_62013 : NOR2A
      port map(A => \General_Controller_0/uc_rx_byte[6]_net_1\, B
         => \General_Controller_0/uc_rx_byte[5]_net_1\, Y => 
        HIEFFPLA_NET_0_74073);
    
    \Science_0/ADC_READ_0/ACLK\ : DFN1E0P1
      port map(D => HIEFFPLA_NET_0_73240, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, E => HIEFFPLA_NET_0_73426, Q => ACLK_c);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/data_out[2]\ : 
        DFN0E1C1
      port map(D => PRESSURE_SDA_in, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72400, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[2]\);
    
    HIEFFPLA_INST_0_63090 : NOR2A
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73831);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[3]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[3]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[3]\);
    
    \Timekeeper_0/microseconds[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72131, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[6]\);
    
    HIEFFPLA_INST_0_59503 : MX2
      port map(A => \Sensors_0_pressure_temp_raw[20]\, B => 
        \Sensors_0_pressure_raw[12]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74545);
    
    \General_Controller_0/st_wen1\ : DFI1E1C1
      port map(D => HIEFFPLA_NET_0_74178, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_74177, CLR => CLKINT_1_Y, QN => 
        \SweepTable_1.WEAP\);
    
    HIEFFPLA_INST_0_55501 : AND2
      port map(A => HIEFFPLA_NET_0_75488, B => 
        HIEFFPLA_NET_0_75486, Y => HIEFFPLA_NET_0_75495);
    
    HIEFFPLA_INST_0_65525 : AND2B
      port map(A => \Science_0/ADC_READ_0/cnt3dn[6]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt3dn[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73352);
    
    HIEFFPLA_INST_0_66981 : OR3A
      port map(A => HIEFFPLA_NET_0_72989, B => 
        HIEFFPLA_NET_0_72974, C => HIEFFPLA_NET_0_72990, Y => 
        HIEFFPLA_NET_0_72991);
    
    HIEFFPLA_INST_0_65364 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt1dn[5]_net_1\, B => 
        HIEFFPLA_NET_0_73413, C => 
        \Science_0/ADC_READ_0/cnt1dn[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73399);
    
    HIEFFPLA_INST_0_57532 : AOI1
      port map(A => \Science_0_exp_packet_0[23]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_75017, Y => HIEFFPLA_NET_0_75018);
    
    \Science_0/DAC_SET_0/state[0]\ : DFN1C1
      port map(D => \Science_0/DAC_SET_0/state[1]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => LDCLK_c);
    
    HIEFFPLA_INST_0_57588 : AOI1
      port map(A => \Science_0_exp_packet_0[43]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74804, Y => HIEFFPLA_NET_0_75000);
    
    \General_Controller_0/sweep_table_samples_per_step[15]\ : 
        DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[15]_net_1\);
    
    HIEFFPLA_INST_0_57138 : AND2
      port map(A => \Sensors_0_pressure_temp_raw[18]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75159);
    
    HIEFFPLA_INST_0_61942 : NOR3B
      port map(A => HIEFFPLA_NET_0_73907, B => 
        HIEFFPLA_NET_0_74073, C => HIEFFPLA_NET_0_73810, Y => 
        HIEFFPLA_NET_0_74092);
    
    \General_Controller_0/readout_en\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74265, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => General_Controller_0_readout_en);
    
    \General_Controller_0/sweep_table_nof_steps[6]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73980, Q => 
        \General_Controller_0/sweep_table_nof_steps[6]_net_1\);
    
    HIEFFPLA_INST_0_57451 : AO1B
      port map(A => \Sensors_0_mag_z[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75041, Y => HIEFFPLA_NET_0_75042);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[3]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72804, Q => 
        \Sensors_0_mag_x[3]\);
    
    HIEFFPLA_INST_0_58023 : AO1
      port map(A => \Science_0_exp_packet_0[73]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75119, Y => HIEFFPLA_NET_0_74876);
    
    HIEFFPLA_INST_0_66081 : AX1
      port map(A => HIEFFPLA_NET_0_73225, B => 
        \Science_0/DAC_SET_0/cnt[3]_net_1\, C => 
        \Science_0/DAC_SET_0/cnt[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73215);
    
    HIEFFPLA_INST_0_69391 : AND3A
      port map(A => HIEFFPLA_NET_0_72429, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        C => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72400);
    
    \Timekeeper_0/microseconds[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72130, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[7]\);
    
    HIEFFPLA_INST_0_59451 : MX2
      port map(A => \Science_0_chan6_data[6]\, B => 
        \Science_0_chan6_data[10]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74553);
    
    HIEFFPLA_INST_0_69620 : AND3B
      port map(A => HIEFFPLA_NET_0_72426, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72343);
    
    HIEFFPLA_INST_0_55036 : NOR3B
      port map(A => HIEFFPLA_NET_0_75600, B => 
        HIEFFPLA_NET_0_75604, C => 
        \Communications_0/UART_0/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75608);
    
    HIEFFPLA_INST_0_66298 : AO1C
      port map(A => HIEFFPLA_NET_0_73166, B => 
        \Science_0/SET_LP_GAIN_0/state[4]_net_1\, C => 
        \Science_0/SET_LP_GAIN_0/state_i_0[0]\, Y => 
        HIEFFPLA_NET_0_73152);
    
    HIEFFPLA_INST_0_70120 : AO1A
      port map(A => HIEFFPLA_NET_0_72271, B => 
        HIEFFPLA_NET_0_72207, C => HIEFFPLA_NET_0_72193, Y => 
        HIEFFPLA_NET_0_72214);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[14]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72283, Q => 
        \Sensors_0_pressure_temp_raw[14]\);
    
    HIEFFPLA_INST_0_69876 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_72239, C => HIEFFPLA_NET_0_72225, Y
         => HIEFFPLA_NET_0_72282);
    
    HIEFFPLA_INST_0_57598 : AOI1
      port map(A => \Science_0_exp_packet_0[44]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74802, Y => HIEFFPLA_NET_0_74997);
    
    HIEFFPLA_INST_0_56559 : AOI1
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/old_acc_new_data_i_0\, B
         => Sensors_0_acc_new_data, C => 
        \Data_Saving_0/Packet_Saver_0/acc_flag_net_1\, Y => 
        HIEFFPLA_NET_0_75239);
    
    HIEFFPLA_INST_0_67362 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\, 
        C => HIEFFPLA_NET_0_72761, Y => HIEFFPLA_NET_0_72898);
    
    HIEFFPLA_INST_0_63728 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[0]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[0]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73721);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[3]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72489, Q => 
        \Sensors_0_gyro_z[3]\);
    
    HIEFFPLA_INST_0_58448 : AOI1
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/old_pressure_new_data_i_0\, 
        B => Sensors_0_pressure_new_data, C => 
        \Data_Saving_0/Packet_Saver_0/pressure_flag_net_1\, Y => 
        HIEFFPLA_NET_0_74764);
    
    HIEFFPLA_INST_0_56474 : XOR3
      port map(A => HIEFFPLA_NET_0_75316, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[0]\\\\\, C => 
        HIEFFPLA_NET_0_75330, Y => HIEFFPLA_NET_0_75271);
    
    HIEFFPLA_INST_0_60708 : MX2
      port map(A => \Science_0_chan5_data[10]\, B => 
        \Science_0_chan4_data[2]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74373);
    
    HIEFFPLA_INST_0_70351 : OR2A
      port map(A => General_Controller_0_st_ren1, B => 
        \SweepTable_0/WEBP\, Y => \SweepTable_1.WEBP\);
    
    HIEFFPLA_INST_0_69609 : AND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        B => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72351);
    
    HIEFFPLA_INST_0_69541 : AO1
      port map(A => 
        \Sensors_0.Pressure_Sensor_0.I2C_Master_0.sda_1\, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_72377, Y => HIEFFPLA_NET_0_72368);
    
    HIEFFPLA_INST_0_67620 : NOR3A
      port map(A => HIEFFPLA_NET_0_72826, B => 
        HIEFFPLA_NET_0_72737, C => HIEFFPLA_NET_0_72736, Y => 
        HIEFFPLA_NET_0_72841);
    
    HIEFFPLA_INST_0_55394 : NAND2B
      port map(A => HIEFFPLA_NET_0_75514, B => 
        HIEFFPLA_NET_0_75527, Y => HIEFFPLA_NET_0_75522);
    
    HIEFFPLA_INST_0_63330 : NOR3A
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        HIEFFPLA_NET_0_73785, C => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73775);
    
    HIEFFPLA_INST_0_69972 : OR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_s_ack_error\, Y
         => HIEFFPLA_NET_0_72256);
    
    HIEFFPLA_INST_0_64656 : NOR3A
      port map(A => HIEFFPLA_NET_0_73606, B => 
        HIEFFPLA_NET_0_73938, C => HIEFFPLA_NET_0_73584, Y => 
        HIEFFPLA_NET_0_73574);
    
    HIEFFPLA_INST_0_60087 : MX2
      port map(A => HIEFFPLA_NET_0_74370, B => 
        HIEFFPLA_NET_0_74398, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74463);
    
    HIEFFPLA_INST_0_70682 : AX1C
      port map(A => HIEFFPLA_NET_0_72038, B => \s_time[5]\, C => 
        \Timing_0/s_time[6]_net_1\, Y => HIEFFPLA_NET_0_72045);
    
    \ClockDivs_0/cnt_800kHz[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75630, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \ClockDivs_0/cnt_800kHz[1]_net_1\);
    
    HIEFFPLA_INST_0_61273 : XA1C
      port map(A => 
        \General_Controller_0/state_seconds[17]_net_1\, B => 
        HIEFFPLA_NET_0_74243, C => HIEFFPLA_NET_0_74217, Y => 
        HIEFFPLA_NET_0_74230);
    
    HIEFFPLA_INST_0_63236 : NAND3C
      port map(A => HIEFFPLA_NET_0_73788, B => 
        \General_Controller_0/uc_rx_substate[4]_net_1\, C => 
        HIEFFPLA_NET_0_73810, Y => HIEFFPLA_NET_0_73801);
    
    \Science_0/ADC_READ_0/cnt1dn[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73403, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1dn[5]_net_1\);
    
    HIEFFPLA_INST_0_61002 : OR3B
      port map(A => \General_Controller_0/ext_rx_state[0]_net_1\, 
        B => \General_Controller_0/ext_rx_state_i_0[1]\, C => 
        Communications_0_ext_rx_rdy, Y => HIEFFPLA_NET_0_74299);
    
    HIEFFPLA_INST_0_55610 : XA1
      port map(A => HIEFFPLA_NET_0_75455, B => 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\, C => 
        HIEFFPLA_NET_0_75437, Y => HIEFFPLA_NET_0_75465);
    
    \General_Controller_0/status_bits_1[61]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74185, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[61]\);
    
    \Data_Saving_0/FPGA_Buffer_0/_RAM4K9_QXI[5]_\ : RAM4K9
      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[7]\\\\\, 
        ADDRA6 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[6]\\\\\, 
        ADDRA5 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\, 
        ADDRA4 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, 
        ADDRA3 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, 
        ADDRA2 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[2]\\\\\, 
        ADDRA1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[1]\\\\\, 
        ADDRA0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[0]\\\\\, 
        ADDRB11 => AFLSDF_GND, ADDRB10 => \GND\, ADDRB9 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\, 
        ADDRB8 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, 
        ADDRB7 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[7]\\\\\, 
        ADDRB6 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, 
        ADDRB5 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\, 
        ADDRB4 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, 
        ADDRB3 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, 
        ADDRB2 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[2]\\\\\, 
        ADDRB1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[1]\\\\\, 
        ADDRB0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[0]\\\\\, 
        DINA8 => \GND\, DINA7 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[29]\, DINA6 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[28]\, DINA5 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[21]\, DINA4 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[20]\, DINA3 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[13]\, DINA2 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[12]\, DINA1 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[5]\, DINA0 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[4]\, DINB8 => 
        \GND\, DINB7 => \GND\, DINB6 => \GND\, DINB5 => \GND\, 
        DINB4 => \GND\, DINB3 => \GND\, DINB2 => \GND\, DINB1 => 
        \GND\, DINB0 => \GND\, WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, 
        WIDTHB0 => \VCC\, WIDTHB1 => \GND\, PIPEA => \GND\, PIPEB
         => \GND\, WMODEA => \GND\, WMODEB => \GND\, BLKA => 
        \Data_Saving_0/FPGA_Buffer_0/MEMWENEG\, BLKB => 
        \AFLSDF_INV_2\, WENA => \GND\, WENB => \VCC\, CLKA => 
        CLKINT_0_Y_0, CLKB => CLKINT_2_Y, RESET => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, DOUTA8 => 
        OPEN, DOUTA7 => OPEN, DOUTA6 => OPEN, DOUTA5 => OPEN, 
        DOUTA4 => OPEN, DOUTA3 => OPEN, DOUTA2 => OPEN, DOUTA1
         => OPEN, DOUTA0 => OPEN, DOUTB8 => OPEN, DOUTB7 => OPEN, 
        DOUTB6 => OPEN, DOUTB5 => OPEN, DOUTB4 => OPEN, DOUTB3
         => OPEN, DOUTB2 => OPEN, DOUTB1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[5]\\\\\, DOUTB0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[4]\\\\\);
    
    HIEFFPLA_INST_0_66705 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_we\, 
        B => HIEFFPLA_NET_0_73049, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73058);
    
    HIEFFPLA_INST_0_55492 : AO1
      port map(A => \Communications_0/UART_0/tx_state[0]_net_1\, 
        B => HIEFFPLA_NET_0_75528, C => HIEFFPLA_NET_0_75497, Y
         => HIEFFPLA_NET_0_75498);
    
    \Data_Saving_0/FPGA_Buffer_0/_RAM4K9_QXI[1]_\ : RAM4K9
      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[7]\\\\\, 
        ADDRA6 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[6]\\\\\, 
        ADDRA5 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\, 
        ADDRA4 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, 
        ADDRA3 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, 
        ADDRA2 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[2]\\\\\, 
        ADDRA1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[1]\\\\\, 
        ADDRA0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[0]\\\\\, 
        ADDRB11 => AFLSDF_GND, ADDRB10 => \GND\, ADDRB9 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\, 
        ADDRB8 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, 
        ADDRB7 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[7]\\\\\, 
        ADDRB6 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, 
        ADDRB5 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\, 
        ADDRB4 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, 
        ADDRB3 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, 
        ADDRB2 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[2]\\\\\, 
        ADDRB1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[1]\\\\\, 
        ADDRB0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[0]\\\\\, 
        DINA8 => \GND\, DINA7 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[25]\, DINA6 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[24]\, DINA5 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[17]\, DINA4 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[16]\, DINA3 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[9]\, DINA2 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[8]\, DINA1 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[1]\, DINA0 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[0]\, DINB8 => 
        \GND\, DINB7 => \GND\, DINB6 => \GND\, DINB5 => \GND\, 
        DINB4 => \GND\, DINB3 => \GND\, DINB2 => \GND\, DINB1 => 
        \GND\, DINB0 => \GND\, WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, 
        WIDTHB0 => \VCC\, WIDTHB1 => \GND\, PIPEA => \GND\, PIPEB
         => \GND\, WMODEA => \GND\, WMODEB => \GND\, BLKA => 
        \Data_Saving_0/FPGA_Buffer_0/MEMWENEG\, BLKB => 
        \AFLSDF_INV_0\, WENA => \GND\, WENB => \VCC\, CLKA => 
        CLKINT_0_Y_0, CLKB => CLKINT_2_Y, RESET => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, DOUTA8 => 
        OPEN, DOUTA7 => OPEN, DOUTA6 => OPEN, DOUTA5 => OPEN, 
        DOUTA4 => OPEN, DOUTA3 => OPEN, DOUTA2 => OPEN, DOUTA1
         => OPEN, DOUTA0 => OPEN, DOUTB8 => OPEN, DOUTB7 => OPEN, 
        DOUTB6 => OPEN, DOUTB5 => OPEN, DOUTB4 => OPEN, DOUTB3
         => OPEN, DOUTB2 => OPEN, DOUTB1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[1]\\\\\, DOUTB0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[0]\\\\\);
    
    HIEFFPLA_INST_0_61100 : AND3C
      port map(A => \Timekeeper_0_milliseconds[13]\, B => 
        \Timekeeper_0_milliseconds[19]\, C => 
        \Timekeeper_0_milliseconds[23]\, Y => 
        HIEFFPLA_NET_0_74277);
    
    \Communications_0/UART_0/rx_rdy\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75551, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75557, Q => 
        \Communications_0/UART_0_rx_rdy\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[14]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72484, Q => 
        \Sensors_0_gyro_y[14]\);
    
    HIEFFPLA_INST_0_69884 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        B => HIEFFPLA_NET_0_72239, C => HIEFFPLA_NET_0_72225, Y
         => HIEFFPLA_NET_0_72280);
    
    HIEFFPLA_INST_0_68809 : NOR3B
      port map(A => HIEFFPLA_NET_0_72477, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, C
         => CLKINT_1_Y, Y => HIEFFPLA_NET_0_72552);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/data_out[1]\ : 
        DFN0E1C1
      port map(D => PRESSURE_SDA_in, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72401, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[1]\);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/temp[7]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72907, Q => 
        \Sensors_0_acc_temp[7]\);
    
    HIEFFPLA_INST_0_66679 : AO1D
      port map(A => HIEFFPLA_NET_0_73047, B => 
        HIEFFPLA_NET_0_73099, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_net_1\, Y
         => HIEFFPLA_NET_0_73067);
    
    HIEFFPLA_INST_0_70791 : AXO7
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_i2c_addr[0]\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72012);
    
    HIEFFPLA_INST_0_62836 : OR3B
      port map(A => HIEFFPLA_NET_0_74113, B => 
        HIEFFPLA_NET_0_74073, C => 
        \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73886);
    
    HIEFFPLA_INST_0_59313 : MX2
      port map(A => \ch3_data_net_0[1]\, B => \ch3_data_net_0[5]\, 
        S => \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74570);
    
    HIEFFPLA_INST_0_70498 : AX1C
      port map(A => \Timekeeper_0_milliseconds[15]\, B => 
        HIEFFPLA_NET_0_72118, C => 
        \Timekeeper_0_milliseconds[16]\, Y => 
        HIEFFPLA_NET_0_72109);
    
    HIEFFPLA_INST_0_66238 : XOR2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G3[0]_net_1\, B
         => \Science_0/ADC_READ_0_G3[0]\, Y => 
        HIEFFPLA_NET_0_73170);
    
    HIEFFPLA_INST_0_59114 : AO1A
      port map(A => HIEFFPLA_NET_0_74382, B => 
        \GS_Readout_0/state[3]_net_1\, C => HIEFFPLA_NET_0_74608, 
        Y => HIEFFPLA_NET_0_74609);
    
    HIEFFPLA_INST_0_65739 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt[3]_net_1\, B => 
        HIEFFPLA_NET_0_73297, C => 
        \Science_0/ADC_READ_0/cnt[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73293);
    
    HIEFFPLA_INST_0_67805 : NOR3A
      port map(A => HIEFFPLA_NET_0_72929, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72797);
    
    HIEFFPLA_INST_0_56378 : AX1D
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, B
         => HIEFFPLA_NET_0_75352, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[7]\\\\\, Y
         => HIEFFPLA_NET_0_75296);
    
    HIEFFPLA_INST_0_70365 : AND3
      port map(A => \Timekeeper_0_microseconds[5]\, B => 
        HIEFFPLA_NET_0_72156, C => \Timekeeper_0_microseconds[6]\, 
        Y => HIEFFPLA_NET_0_72159);
    
    HIEFFPLA_INST_0_59285 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[41]\, B => 
        \Data_Hub_Packets_0_status_packet[45]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74575);
    
    HIEFFPLA_INST_0_63946 : MX2
      port map(A => HIEFFPLA_NET_0_73657, B => 
        HIEFFPLA_NET_0_73649, S => HIEFFPLA_NET_0_73599, Y => 
        HIEFFPLA_NET_0_73686);
    
    HIEFFPLA_INST_0_61041 : AO1A
      port map(A => \General_Controller_0/mission_mode_net_1\, B
         => \General_Controller_0/flight_state[3]_net_1\, C => 
        HIEFFPLA_NET_0_74288, Y => HIEFFPLA_NET_0_74289);
    
    HIEFFPLA_INST_0_68379 : OR2A
      port map(A => HIEFFPLA_NET_0_72689, B => GYRO_SCL_c, Y => 
        HIEFFPLA_NET_0_72664);
    
    HIEFFPLA_INST_0_55699 : AND2B
      port map(A => \Communications_0/UART_1/rx_state[0]_net_1\, 
        B => \Communications_0/UART_1/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75443);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[7]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72808, Q => 
        \Sensors_0_mag_z[7]\);
    
    HIEFFPLA_INST_0_66086 : NAND2B
      port map(A => \Science_0/DAC_SET_0/state[1]_net_1\, B => 
        HIEFFPLA_NET_0_73226, Y => HIEFFPLA_NET_0_73212);
    
    HIEFFPLA_INST_0_62932 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => \General_Controller_0/uc_rx_substate[2]_net_1\, C
         => HIEFFPLA_NET_0_73810, Y => HIEFFPLA_NET_0_73864);
    
    \General_Controller_0/sweep_table_write_value[13]\ : DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[13]_net_1\);
    
    \Science_0/ADC_READ_0/cnt2up[0]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73364, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2up[0]_net_1\);
    
    \General_Controller_0/sweep_table_sweep_cnt[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74133, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[5]_net_1\);
    
    \AA_pad/U0/U1\ : IOIN_IB
      port map(YIN => \AA_pad/U0/NET1\, Y => AA_c);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[6]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[6]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[6]\);
    
    HIEFFPLA_INST_0_66650 : OR3B
      port map(A => HIEFFPLA_NET_0_73045, B => 
        HIEFFPLA_NET_0_73042, C => HIEFFPLA_NET_0_73072, Y => 
        HIEFFPLA_NET_0_73073);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72333, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\);
    
    HIEFFPLA_INST_0_64829 : AX1B
      port map(A => HIEFFPLA_NET_0_73523, B => 
        HIEFFPLA_NET_0_73526, C => 
        \General_Controller_0/uc_tx_substate[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73529);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[0]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[0]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[0]\);
    
    HIEFFPLA_INST_0_70714 : AND2
      port map(A => \Timing_0/s_time[2]_net_1\, B => 
        \s_clks_net_0[18]\, Y => HIEFFPLA_NET_0_72034);
    
    HIEFFPLA_INST_0_65130 : NAND2B
      port map(A => \Sensors_0_pressure_raw[20]\, B => 
        \Sensors_0_pressure_raw[21]\, Y => HIEFFPLA_NET_0_73463);
    
    HIEFFPLA_INST_0_69859 : AOI1C
      port map(A => \Sensors_0/Pressure_Sensor_0/state[8]\, B => 
        HIEFFPLA_NET_0_72244, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        Y => HIEFFPLA_NET_0_72288);
    
    \GS_Readout_0/prevState[0]\ : DFN1E0C1
      port map(D => \GS_Readout_0/state[0]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \GS_Readout_0/state[6]_net_1\, Q => 
        \GS_Readout_0/prevState[0]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/num_bytes_1[2]\ : 
        DFN1
      port map(D => HIEFFPLA_NET_0_72965, CLK => CLKINT_0_Y_0, Q
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[2]\);
    
    HIEFFPLA_INST_0_69017 : NAND3A
      port map(A => CLKINT_1_Y, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        C => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72497);
    
    HIEFFPLA_INST_0_57815 : NAND3C
      port map(A => HIEFFPLA_NET_0_74825, B => 
        HIEFFPLA_NET_0_74809, C => HIEFFPLA_NET_0_74776, Y => 
        HIEFFPLA_NET_0_74935);
    
    HIEFFPLA_INST_0_70668 : XA1B
      port map(A => HIEFFPLA_NET_0_72022, B => 
        \Timing_0/s_count[7]_net_1\, C => HIEFFPLA_NET_0_72058, Y
         => HIEFFPLA_NET_0_72050);
    
    HIEFFPLA_INST_0_68356 : AND3A
      port map(A => HIEFFPLA_NET_0_72703, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, C => 
        GYRO_SCL_c, Y => HIEFFPLA_NET_0_72673);
    
    HIEFFPLA_INST_0_62492 : NOR3B
      port map(A => HIEFFPLA_NET_0_73888, B => 
        HIEFFPLA_NET_0_73906, C => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73971);
    
    \LA1_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => LA1_c, E => \VCC\, DOUT => \LA1_pad/U0/NET1\, 
        EOUT => \LA1_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_57161 : AND2
      port map(A => \ch3_data_net_0[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75144);
    
    HIEFFPLA_INST_0_69971 : OR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[3]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_s_ack_error\, Y
         => HIEFFPLA_NET_0_72257);
    
    HIEFFPLA_INST_0_58350 : AO1
      port map(A => \Sensors_0_mag_x[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75086, Y => HIEFFPLA_NET_0_74795);
    
    HIEFFPLA_INST_0_67013 : AOI1D
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, B
         => HIEFFPLA_NET_0_72884, C => HIEFFPLA_NET_0_72977, Y
         => HIEFFPLA_NET_0_72985);
    
    HIEFFPLA_INST_0_58599 : AX1B
      port map(A => \GS_Readout_0/subState[3]_net_1\, B => 
        HIEFFPLA_NET_0_74343, C => 
        \GS_Readout_0/subState[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74725);
    
    HIEFFPLA_INST_0_56968 : MX2
      port map(A => HIEFFPLA_NET_0_74967, B => 
        HIEFFPLA_NET_0_74897, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75189);
    
    HIEFFPLA_INST_0_63614 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[13]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_sample_skip[13]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73740);
    
    HIEFFPLA_INST_0_63009 : AND3
      port map(A => HIEFFPLA_NET_0_74070, B => 
        \General_Controller_0/uc_rx_state_0[1]_net_1\, C => 
        HIEFFPLA_NET_0_74026, Y => HIEFFPLA_NET_0_73848);
    
    \Science_0/SET_LP_GAIN_0/old_G3[0]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73169, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/old_G3[0]_net_1\);
    
    \Science_0/ADC_READ_0/chan4_data[2]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[2]\);
    
    HIEFFPLA_INST_0_62361 : NAND3C
      port map(A => HIEFFPLA_NET_0_73942, B => 
        HIEFFPLA_NET_0_74096, C => HIEFFPLA_NET_0_73976, Y => 
        HIEFFPLA_NET_0_73997);
    
    \FFU_EJECTED_pad/U0/U1\ : IOIN_IB
      port map(YIN => \FFU_EJECTED_pad/U0/NET1\, Y => 
        FFU_EJECTED_c);
    
    HIEFFPLA_INST_0_67184 : AND3
      port map(A => HIEFFPLA_NET_0_72954, B => 
        HIEFFPLA_NET_0_72958, C => HIEFFPLA_NET_0_72950, Y => 
        HIEFFPLA_NET_0_72944);
    
    HIEFFPLA_INST_0_55459 : XA1B
      port map(A => \Communications_0/UART_0/tx_count[0]_net_1\, 
        B => \Communications_0/UART_0/tx_count[1]_net_1\, C => 
        HIEFFPLA_NET_0_75502, Y => HIEFFPLA_NET_0_75506);
    
    HIEFFPLA_INST_0_63656 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[12]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_samples_per_point[12]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73733);
    
    HIEFFPLA_INST_0_59081 : AND3
      port map(A => HIEFFPLA_NET_0_74615, B => 
        HIEFFPLA_NET_0_74510, C => HIEFFPLA_NET_0_74435, Y => 
        HIEFFPLA_NET_0_74618);
    
    HIEFFPLA_INST_0_66736 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        B => HIEFFPLA_NET_0_73101, Y => HIEFFPLA_NET_0_73050);
    
    HIEFFPLA_INST_0_63476 : MX2
      port map(A => HIEFFPLA_NET_0_73684, B => 
        HIEFFPLA_NET_0_73676, S => HIEFFPLA_NET_0_73621, Y => 
        HIEFFPLA_NET_0_73759);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/write_done\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72422, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72318, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_write_done\);
    
    HIEFFPLA_INST_0_65651 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt4dn[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt4dn[0]_net_1\, C => 
        HIEFFPLA_NET_0_73274, Y => HIEFFPLA_NET_0_73317);
    
    HIEFFPLA_INST_0_63286 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state_0[1]_net_1\, 
        B => HIEFFPLA_NET_0_73897, C => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73787);
    
    HIEFFPLA_INST_0_62025 : NOR3B
      port map(A => HIEFFPLA_NET_0_74069, B => 
        HIEFFPLA_NET_0_73882, C => HIEFFPLA_NET_0_73889, Y => 
        HIEFFPLA_NET_0_74068);
    
    HIEFFPLA_INST_0_55367 : AO1
      port map(A => HIEFFPLA_NET_0_75531, B => 
        HIEFFPLA_NET_0_75530, C => 
        \Communications_0/UART_0/tx_clk_count_i_0[8]\, Y => 
        HIEFFPLA_NET_0_75528);
    
    HIEFFPLA_INST_0_66747 : MX2
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_73044, S => ACCE_SCL_c, Y => 
        HIEFFPLA_NET_0_73047);
    
    HIEFFPLA_INST_0_57802 : AO1
      port map(A => \Sensors_0_gyro_x[15]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74937, Y => HIEFFPLA_NET_0_74938);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[0]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72489, Q => 
        \Sensors_0_gyro_z[0]\);
    
    HIEFFPLA_INST_0_60865 : AND2
      port map(A => HIEFFPLA_NET_0_74333, B => 
        HIEFFPLA_NET_0_74326, Y => HIEFFPLA_NET_0_74336);
    
    HIEFFPLA_INST_0_68890 : NOR3B
      port map(A => HIEFFPLA_NET_0_72508, B => 
        HIEFFPLA_NET_0_72530, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72531);
    
    HIEFFPLA_INST_0_70319 : AO1A
      port map(A => HIEFFPLA_NET_0_72278, B => 
        HIEFFPLA_NET_0_72188, C => HIEFFPLA_NET_0_72174, Y => 
        HIEFFPLA_NET_0_72175);
    
    \Eject_Signal_Debounce_0/state[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74735, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72220, Q => 
        \Eject_Signal_Debounce_0/state[0]_net_1\);
    
    HIEFFPLA_INST_0_70024 : AO1C
      port map(A => HIEFFPLA_NET_0_72284, B => 
        HIEFFPLA_NET_0_72285, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72244);
    
    HIEFFPLA_INST_0_57986 : AO1
      port map(A => \Science_0_exp_packet_0[31]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74784, Y => HIEFFPLA_NET_0_74887);
    
    HIEFFPLA_INST_0_57631 : AO1B
      port map(A => \Sensors_0_acc_y[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74986, Y => HIEFFPLA_NET_0_74987);
    
    HIEFFPLA_INST_0_55717 : AO1A
      port map(A => \Communications_0/UART_1/rx_state[0]_net_1\, 
        B => HIEFFPLA_NET_0_75482, C => HIEFFPLA_NET_0_75439, Y
         => HIEFFPLA_NET_0_75438);
    
    HIEFFPLA_INST_0_71014 : XA1C
      port map(A => Communications_0_uc_tx_rdy, B => 
        \General_Controller_0/uc_tx_substate[0]_net_1\, C => 
        HIEFFPLA_NET_0_71988, Y => HIEFFPLA_NET_0_73542);
    
    HIEFFPLA_INST_0_70968 : MX2A
      port map(A => HIEFFPLA_NET_0_71999, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[2]\, 
        S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_73128);
    
    HIEFFPLA_INST_0_65527 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt3dn[4]_net_1\, B => 
        HIEFFPLA_NET_0_73348, C => 
        \Science_0/ADC_READ_0/cnt3dn[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73351);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/data_out_1[2]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_72568, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72547, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[2]\);
    
    HIEFFPLA_INST_0_65487 : NOR3A
      port map(A => HIEFFPLA_NET_0_73276, B => 
        \Science_0/ADC_READ_0/cnt2up[0]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt2up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73364);
    
    HIEFFPLA_INST_0_62375 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        HIEFFPLA_NET_0_73889, Y => HIEFFPLA_NET_0_73994);
    
    \UC_UART_TX_pad/U0/U1\ : IOIN_IB
      port map(YIN => \UC_UART_TX_pad/U0/NET1\, Y => UC_UART_TX_c);
    
    HIEFFPLA_INST_0_71062 : NAND3C
      port map(A => \General_Controller_0/state_seconds[2]_net_1\, 
        B => \General_Controller_0/state_seconds[1]_net_1\, C => 
        \General_Controller_0/state_seconds[8]_net_1\, Y => 
        HIEFFPLA_NET_0_71984);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRY[5]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75289, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[5]\\\\\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[3]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[3]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[3]\);
    
    HIEFFPLA_INST_0_55999 : NAND3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, B
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\, 
        C => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, 
        Y => HIEFFPLA_NET_0_75373);
    
    HIEFFPLA_INST_0_88379 : MIN3
      port map(A => HIEFFPLA_NET_0_75288, B => 
        HIEFFPLA_NET_0_75321, C => HIEFFPLA_NET_0_89694, Y => 
        HIEFFPLA_NET_0_88380);
    
    HIEFFPLA_INST_0_55909 : NAND2B
      port map(A => HIEFFPLA_NET_0_75414, B => 
        \Communications_0/UART_1/tx_clk_count_i_0[7]\, Y => 
        HIEFFPLA_NET_0_75398);
    
    HIEFFPLA_INST_0_63776 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[0]_net_1\, 
        B => \General_Controller_0/sweep_table_points[0]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73713);
    
    HIEFFPLA_INST_0_62244 : AOI1
      port map(A => HIEFFPLA_NET_0_73793, B => 
        HIEFFPLA_NET_0_73909, C => HIEFFPLA_NET_0_74021, Y => 
        HIEFFPLA_NET_0_74022);
    
    HIEFFPLA_INST_0_69622 : NAND3C
      port map(A => HIEFFPLA_NET_0_72343, B => 
        HIEFFPLA_NET_0_72344, C => HIEFFPLA_NET_0_72425, Y => 
        HIEFFPLA_NET_0_72342);
    
    HIEFFPLA_INST_0_61085 : OR3B
      port map(A => HIEFFPLA_NET_0_74275, B => 
        HIEFFPLA_NET_0_74280, C => 
        \Timekeeper_0_milliseconds[11]\, Y => 
        HIEFFPLA_NET_0_74281);
    
    HIEFFPLA_INST_0_62031 : NAND3C
      port map(A => HIEFFPLA_NET_0_73858, B => 
        HIEFFPLA_NET_0_73859, C => HIEFFPLA_NET_0_74066, Y => 
        HIEFFPLA_NET_0_74067);
    
    HIEFFPLA_INST_0_58404 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[40]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_74777);
    
    HIEFFPLA_INST_0_57082 : MX2
      port map(A => HIEFFPLA_NET_0_74941, B => CU_SYNC_c, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75171);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/isSetup\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72313, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/isSetup_net_1\);
    
    HIEFFPLA_INST_0_70793 : MX2
      port map(A => HIEFFPLA_NET_0_72370, B => 
        HIEFFPLA_NET_0_72367, S => PRESSURE_SCL_c, Y => 
        HIEFFPLA_NET_0_72011);
    
    HIEFFPLA_INST_0_67676 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72826);
    
    HIEFFPLA_INST_0_67153 : AND3C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72950);
    
    HIEFFPLA_INST_0_67895 : OA1C
      port map(A => HIEFFPLA_NET_0_72743, B => 
        HIEFFPLA_NET_0_72792, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, Y
         => HIEFFPLA_NET_0_72778);
    
    HIEFFPLA_INST_0_59236 : AND2
      port map(A => \GS_Readout_0/state[0]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74582);
    
    HIEFFPLA_INST_0_68562 : AO1D
      port map(A => HIEFFPLA_NET_0_72698, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, C => 
        HIEFFPLA_NET_0_72628, Y => HIEFFPLA_NET_0_72617);
    
    HIEFFPLA_INST_0_62169 : NOR3A
      port map(A => HIEFFPLA_NET_0_73993, B => 
        HIEFFPLA_NET_0_74042, C => HIEFFPLA_NET_0_74037, Y => 
        HIEFFPLA_NET_0_74038);
    
    \GS_Readout_0/subState[0]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_74356, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => \GS_Readout_0/subState_0[0]\);
    
    HIEFFPLA_INST_0_66912 : NAND3B
      port map(A => HIEFFPLA_NET_0_72793, B => 
        HIEFFPLA_NET_0_72750, C => HIEFFPLA_NET_0_72911, Y => 
        HIEFFPLA_NET_0_73006);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[11]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72782, Q => 
        \Sensors_0_mag_y[11]\);
    
    HIEFFPLA_INST_0_68690 : NAND2B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72586);
    
    HIEFFPLA_INST_0_69435 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[2]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72390);
    
    HIEFFPLA_INST_0_69153 : NOR3A
      port map(A => \Sensors_0/Gyro_0/state[8]\, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        C => HIEFFPLA_NET_0_72540, Y => HIEFFPLA_NET_0_72459);
    
    HIEFFPLA_INST_0_65579 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt3dn[6]_net_1\, B => 
        HIEFFPLA_NET_0_73351, C => 
        \Science_0/ADC_READ_0/cnt3dn[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73339);
    
    \ClockDivs_0/clk_800kHz\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75637, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \ClockDivs_0/clk_800kHz_i\);
    
    HIEFFPLA_INST_0_62743 : XOR2
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73916);
    
    HIEFFPLA_INST_0_59030 : AO1A
      port map(A => HIEFFPLA_NET_0_74552, B => 
        HIEFFPLA_NET_0_74660, C => HIEFFPLA_NET_0_74631, Y => 
        HIEFFPLA_NET_0_74632);
    
    HIEFFPLA_INST_0_68087 : AND2
      port map(A => HIEFFPLA_NET_0_72886, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, Y
         => HIEFFPLA_NET_0_72732);
    
    HIEFFPLA_INST_0_54962 : AO1E
      port map(A => 
        \Communications_0/FFU_Command_Checker_0/state[0]_net_1\, 
        B => \Communications_0/UART_0_rx_rdy\, C => 
        \Communications_0/FFU_Command_Checker_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_75626);
    
    \Science_0/ADC_READ_0/chan[1]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/cnt_chan[1]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73238, Q => 
        \Science_0/ADC_READ_0/chan[1]_net_1\);
    
    \Science_0/DAC_SET_0/state[1]\ : DFN1C1
      port map(D => \Science_0/DAC_SET_0/state[2]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_68080 : XAI1
      port map(A => HIEFFPLA_NET_0_72921, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        C => HIEFFPLA_NET_0_72758, Y => HIEFFPLA_NET_0_72735);
    
    HIEFFPLA_INST_0_70440 : XOR2
      port map(A => HIEFFPLA_NET_0_72157, B => 
        \Timekeeper_0_microseconds[9]\, Y => HIEFFPLA_NET_0_72128);
    
    HIEFFPLA_INST_0_61855 : AXOI3
      port map(A => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_byte[3]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74115);
    
    \Data_Saving_0/Packet_Saver_0/data_out[4]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75209, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[4]\);
    
    HIEFFPLA_INST_0_68323 : AND3C
      port map(A => HIEFFPLA_NET_0_72676, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72682);
    
    HIEFFPLA_INST_0_57454 : AOI1
      port map(A => \Science_0_exp_packet_0[27]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_75040, Y => HIEFFPLA_NET_0_75041);
    
    HIEFFPLA_INST_0_69076 : NOR3A
      port map(A => HIEFFPLA_NET_0_72540, B => CLKINT_1_Y, C => 
        HIEFFPLA_NET_0_72488, Y => HIEFFPLA_NET_0_72476);
    
    \Communications_0/UART_0/tx_count[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75507, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75503, Q => 
        \Communications_0/UART_0/tx_count[1]_net_1\);
    
    HIEFFPLA_INST_0_58947 : NAND3C
      port map(A => HIEFFPLA_NET_0_74645, B => 
        HIEFFPLA_NET_0_74484, C => HIEFFPLA_NET_0_74646, Y => 
        HIEFFPLA_NET_0_74651);
    
    HIEFFPLA_INST_0_56490 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[1]\\\\\, B
         => HIEFFPLA_NET_0_75369, Y => HIEFFPLA_NET_0_75266);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[7]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72489, Q => 
        \ch3_data_net_0[3]\);
    
    \LED2_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => LED2_c, E => \VCC\, DOUT => 
        \LED2_pad/U0/NET1\, EOUT => \LED2_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_67482 : AO1A
      port map(A => HIEFFPLA_NET_0_72853, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        C => HIEFFPLA_NET_0_72867, Y => HIEFFPLA_NET_0_72868);
    
    HIEFFPLA_INST_0_59454 : NOR2A
      port map(A => HIEFFPLA_NET_0_74472, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74552);
    
    \General_Controller_0/uc_rx_byte[3]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[3]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte[3]_net_1\);
    
    HIEFFPLA_INST_0_59985 : MX2
      port map(A => \ch3_data_net_0[9]\, B => 
        \Sensors_0_acc_z[1]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74478);
    
    \General_Controller_0/sweep_table_samples_per_point[6]\ : 
        DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[6]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[6]_net_1\);
    
    \General_Controller_0/uc_tx_state[12]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73574, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[12]_net_1\);
    
    HIEFFPLA_INST_0_58029 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_74873);
    
    \General_Controller_0/status_bits_1[52]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74194, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[52]\);
    
    \Communications_0/UART_1/tx_byte[1]\ : DFN1E1
      port map(D => \General_Controller_0_uc_send[1]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_75385, Q => 
        \Communications_0/UART_1/tx_byte[1]_net_1\);
    
    HIEFFPLA_INST_0_62617 : OR2A
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => Communications_0_uc_rx_rdy, Y => 
        HIEFFPLA_NET_0_73944);
    
    HIEFFPLA_INST_0_60470 : MX2
      port map(A => HIEFFPLA_NET_0_74475, B => 
        HIEFFPLA_NET_0_74463, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74410);
    
    HIEFFPLA_INST_0_56982 : AOI1D
      port map(A => HIEFFPLA_NET_0_74845, B => 
        HIEFFPLA_NET_0_74962, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75187);
    
    \Science_0/ADC_READ_0/chan[0]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/cnt_chan[0]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73238, Q => 
        \Science_0/ADC_READ_0/chan[0]_net_1\);
    
    HIEFFPLA_INST_0_70404 : AX1C
      port map(A => \Timekeeper_0_microseconds[13]\, B => 
        HIEFFPLA_NET_0_72155, C => 
        \Timekeeper_0_microseconds[14]\, Y => 
        HIEFFPLA_NET_0_72146);
    
    HIEFFPLA_INST_0_68438 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[5]_net_1\, B => 
        HIEFFPLA_NET_0_72700, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, Y => 
        HIEFFPLA_NET_0_72650);
    
    \Science_0/ADC_READ_0/exp_packet_1[31]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[15]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[31]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[11]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72553, Q => 
        \Sensors_0_gyro_x[11]\);
    
    HIEFFPLA_INST_0_65483 : NAND3
      port map(A => HIEFFPLA_NET_0_73276, B => 
        \Science_0/ADC_READ_0/cnt2up[4]_net_1\, C => 
        \Science_0/ADC_READ_0_G2[0]\, Y => HIEFFPLA_NET_0_73365);
    
    HIEFFPLA_INST_0_68843 : NOR3B
      port map(A => HIEFFPLA_NET_0_72541, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, C
         => CLKINT_1_Y, Y => HIEFFPLA_NET_0_72542);
    
    HIEFFPLA_INST_0_68633 : AND3C
      port map(A => HIEFFPLA_NET_0_72705, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_72601);
    
    HIEFFPLA_INST_0_59136 : NOR3B
      port map(A => HIEFFPLA_NET_0_74719, B => 
        \GS_Readout_0/prevState[4]_net_1\, C => 
        \GS_Readout_0/prevState[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74603);
    
    \General_Controller_0/st_wdata[6]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[6]\);
    
    HIEFFPLA_INST_0_54965 : NOR3B
      port map(A => 
        \Communications_0/FFU_Command_Checker_0/state[1]_net_1\, 
        B => \Communications_0/UART_0_rx_rdy\, C => 
        \Communications_0/FFU_Command_Checker_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_75625);
    
    HIEFFPLA_INST_0_55791 : MX2
      port map(A => HIEFFPLA_NET_0_75422, B => 
        HIEFFPLA_NET_0_75421, S => 
        \Communications_0/UART_1/tx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75425);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_72418, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\);
    
    HIEFFPLA_INST_0_63506 : MX2
      port map(A => HIEFFPLA_NET_0_73681, B => 
        HIEFFPLA_NET_0_73673, S => HIEFFPLA_NET_0_73621, Y => 
        HIEFFPLA_NET_0_73756);
    
    HIEFFPLA_INST_0_57809 : NAND3C
      port map(A => HIEFFPLA_NET_0_74827, B => 
        HIEFFPLA_NET_0_74810, C => HIEFFPLA_NET_0_74778, Y => 
        HIEFFPLA_NET_0_74936);
    
    \General_Controller_0/sweep_table_write_wait[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74123, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/sweep_table_write_wait[0]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRYSYNC[0]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_10_Q\, 
        CLK => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[0]\\\\\);
    
    HIEFFPLA_INST_0_63182 : NOR3B
      port map(A => HIEFFPLA_NET_0_73779, B => 
        HIEFFPLA_NET_0_73918, C => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_73814);
    
    HIEFFPLA_INST_0_60905 : OR3A
      port map(A => HIEFFPLA_NET_0_74319, B => 
        \General_Controller_0/un10_uc_tx_rdy_i[3]\, C => 
        \General_Controller_0/un10_uc_tx_rdy_i[2]\, Y => 
        HIEFFPLA_NET_0_74323);
    
    HIEFFPLA_INST_0_69581 : AND3C
      port map(A => HIEFFPLA_NET_0_72358, B => 
        HIEFFPLA_NET_0_72357, C => HIEFFPLA_NET_0_72425, Y => 
        HIEFFPLA_NET_0_72359);
    
    HIEFFPLA_INST_0_55931 : AO1A
      port map(A => HIEFFPLA_NET_0_75387, B => 
        HIEFFPLA_NET_0_75389, C => HIEFFPLA_NET_0_75396, Y => 
        HIEFFPLA_NET_0_75392);
    
    HIEFFPLA_INST_0_61452 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[49]\, B => 
        \Timekeeper_0_milliseconds[9]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74197);
    
    HIEFFPLA_INST_0_63354 : MX2A
      port map(A => HIEFFPLA_NET_0_74000, B => 
        HIEFFPLA_NET_0_73536, S => HIEFFPLA_NET_0_73965, Y => 
        HIEFFPLA_NET_0_73772);
    
    HIEFFPLA_INST_0_65560 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt3dn[4]_net_1\, B => 
        HIEFFPLA_NET_0_73357, C => HIEFFPLA_NET_0_73349, Y => 
        HIEFFPLA_NET_0_73343);
    
    HIEFFPLA_INST_0_63197 : OR2A
      port map(A => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73811);
    
    HIEFFPLA_INST_0_59275 : MX2
      port map(A => HIEFFPLA_NET_0_74561, B => 
        HIEFFPLA_NET_0_74551, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74576);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_new_data\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72968, Q => Sensors_0_mag_new_data);
    
    HIEFFPLA_INST_0_66259 : MX2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G4[0]_net_1\, B
         => \Science_0/ADC_READ_0_G4[0]\, S => 
        \Science_0/SET_LP_GAIN_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73164);
    
    HIEFFPLA_INST_0_66375 : OR3A
      port map(A => HIEFFPLA_NET_0_73134, B => 
        HIEFFPLA_NET_0_73039, C => HIEFFPLA_NET_0_73133, Y => 
        HIEFFPLA_NET_0_73135);
    
    HIEFFPLA_INST_0_57372 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_74853, Y => HIEFFPLA_NET_0_75064);
    
    HIEFFPLA_INST_0_59141 : NOR3B
      port map(A => HIEFFPLA_NET_0_74591, B => 
        \GS_Readout_0/subState[1]_net_1\, C => 
        \GS_Readout_0/subState[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74602);
    
    HIEFFPLA_INST_0_56430 : MX2
      port map(A => \FMC_DA_c[4]\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[4]\\\\\, S => 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\, Y => 
        HIEFFPLA_NET_0_75283);
    
    HIEFFPLA_INST_0_67908 : OR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72775);
    
    HIEFFPLA_INST_0_56339 : AX1D
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\, B
         => HIEFFPLA_NET_0_75257, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[10]\\\\\, Y
         => HIEFFPLA_NET_0_75306);
    
    HIEFFPLA_INST_0_61292 : AOI1D
      port map(A => HIEFFPLA_NET_0_74295, B => 
        HIEFFPLA_NET_0_74293, C => HIEFFPLA_NET_0_74214, Y => 
        HIEFFPLA_NET_0_74226);
    
    HIEFFPLA_INST_0_59838 : OA1C
      port map(A => HIEFFPLA_NET_0_74433, B => 
        HIEFFPLA_NET_0_74725, C => HIEFFPLA_NET_0_74574, Y => 
        HIEFFPLA_NET_0_74500);
    
    HIEFFPLA_INST_0_67414 : NOR3A
      port map(A => HIEFFPLA_NET_0_72889, B => 
        HIEFFPLA_NET_0_72739, C => HIEFFPLA_NET_0_72799, Y => 
        HIEFFPLA_NET_0_72887);
    
    HIEFFPLA_INST_0_61311 : XA1B
      port map(A => \General_Controller_0/state_seconds[6]_net_1\, 
        B => HIEFFPLA_NET_0_74212, C => HIEFFPLA_NET_0_74217, Y
         => HIEFFPLA_NET_0_74221);
    
    HIEFFPLA_INST_0_70066 : AO1C
      port map(A => HIEFFPLA_NET_0_72311, B => 
        HIEFFPLA_NET_0_72302, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        Y => HIEFFPLA_NET_0_72230);
    
    HIEFFPLA_INST_0_60049 : AND2
      port map(A => HIEFFPLA_NET_0_74474, B => 
        HIEFFPLA_NET_0_74552, Y => HIEFFPLA_NET_0_74469);
    
    HIEFFPLA_INST_0_57093 : AOI1C
      port map(A => HIEFFPLA_NET_0_74938, B => 
        HIEFFPLA_NET_0_74883, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75168);
    
    HIEFFPLA_INST_0_70635 : AND3A
      port map(A => HIEFFPLA_NET_0_72060, B => 
        \Timing_0/s_count[5]_net_1\, C => 
        \Timing_0/s_count[4]_net_1\, Y => HIEFFPLA_NET_0_72057);
    
    HIEFFPLA_INST_0_65586 : AND2
      port map(A => \Science_0/ADC_READ_0/cnt3up[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt3up[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73337);
    
    HIEFFPLA_INST_0_56937 : MX2
      port map(A => HIEFFPLA_NET_0_74978, B => 
        HIEFFPLA_NET_0_74906, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75193);
    
    \General_Controller_0/command[6]\ : DFN1E1
      port map(D => \Communications_0_ext_recv[6]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74300, Q => 
        \General_Controller_0/command[6]_net_1\);
    
    HIEFFPLA_INST_0_67065 : NAND2B
      port map(A => \Sensors_0/Accelerometer_0/state_0[8]\, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[3]\, 
        Y => HIEFFPLA_NET_0_72973);
    
    \Science_0/SET_LP_GAIN_0/LA0\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_73185, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73160, Q => LA0_c);
    
    HIEFFPLA_INST_0_64112 : OR2A
      port map(A => HIEFFPLA_NET_0_73579, B => 
        \General_Controller_0/constant_bias_voltage_0[12]_net_1\, 
        Y => HIEFFPLA_NET_0_73668);
    
    HIEFFPLA_INST_0_70227 : AO1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_write_done\, C
         => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72191);
    
    HIEFFPLA_INST_0_65291 : NAND3
      port map(A => \Science_0/ADC_READ_0/newflag_net_1\, B => 
        \Science_0/ADC_READ_0/chan[0]_net_1\, C => 
        \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73421);
    
    HIEFFPLA_INST_0_63121 : AND3
      port map(A => HIEFFPLA_NET_0_73823, B => 
        HIEFFPLA_NET_0_74092, C => HIEFFPLA_NET_0_74026, Y => 
        HIEFFPLA_NET_0_73824);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[16]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[16]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[16]\);
    
    HIEFFPLA_INST_0_62885 : OR3A
      port map(A => \General_Controller_0/uc_rx_state[1]_net_1\, 
        B => \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73875);
    
    HIEFFPLA_INST_0_56528 : XOR2
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[0]_net_1\, B
         => 
        \Data_Saving_0/Interrupt_Generator_0/counter[1]_net_1\, Y
         => HIEFFPLA_NET_0_75252);
    
    \Science_0/ADC_READ_0/chan1_data[7]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[7]\);
    
    \General_Controller_0/temp_first_byte[6]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73872, Q => 
        \General_Controller_0/temp_first_byte[6]_net_1\);
    
    HIEFFPLA_INST_0_71217 : AXOI1
      port map(A => HIEFFPLA_NET_0_75619, B => 
        HIEFFPLA_NET_0_71971, C => HIEFFPLA_NET_0_71970, Y => 
        HIEFFPLA_NET_0_75623);
    
    HIEFFPLA_INST_0_69890 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[1]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72278);
    
    HIEFFPLA_INST_0_62834 : NOR2A
      port map(A => \General_Controller_0/uc_rx_state[3]_net_1\, 
        B => \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73887);
    
    \Sensors_0/Gyro_0/I2C_Master_0/state[2]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72611, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[2]_net_1\);
    
    HIEFFPLA_INST_0_61208 : AND2
      port map(A => 
        \General_Controller_0/state_seconds[15]_net_1\, B => 
        \General_Controller_0/state_seconds[14]_net_1\, Y => 
        HIEFFPLA_NET_0_74250);
    
    \Science_0/ADC_READ_0/cnt4up[3]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73302, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4up[3]_net_1\);
    
    HIEFFPLA_INST_0_55571 : AND3C
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[26]_net_1\, B => 
        \Communications_0/UART_1/rx_clk_count[27]_net_1\, C => 
        \Communications_0/UART_1/rx_clk_count[25]_net_1\, Y => 
        HIEFFPLA_NET_0_75478);
    
    HIEFFPLA_INST_0_69517 : AND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72373);
    
    \General_Controller_0/st_waddr[5]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[5]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_waddr[5]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[78]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[22]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[78]\);
    
    HIEFFPLA_INST_0_59071 : NOR3B
      port map(A => HIEFFPLA_NET_0_74521, B => 
        HIEFFPLA_NET_0_74510, C => HIEFFPLA_NET_0_74450, Y => 
        HIEFFPLA_NET_0_74622);
    
    \Science_0/ADC_READ_0/cnt2dn[3]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73373, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2dn[3]_net_1\);
    
    HIEFFPLA_INST_0_61428 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[46]\, B => 
        \Timekeeper_0_milliseconds[6]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74200);
    
    HIEFFPLA_INST_0_70521 : AX1C
      port map(A => \Timekeeper_0_milliseconds[3]\, B => 
        HIEFFPLA_NET_0_72125, C => \Timekeeper_0_milliseconds[4]\, 
        Y => HIEFFPLA_NET_0_72098);
    
    HIEFFPLA_INST_0_65453 : XA1C
      port map(A => \Science_0/ADC_READ_0/cnt2dn[4]_net_1\, B => 
        HIEFFPLA_NET_0_73387, C => HIEFFPLA_NET_0_73381, Y => 
        HIEFFPLA_NET_0_73372);
    
    HIEFFPLA_INST_0_56095 : NOR3B
      port map(A => HIEFFPLA_NET_0_75376, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, C
         => HIEFFPLA_NET_0_75370, Y => HIEFFPLA_NET_0_75348);
    
    \Science_0/ADC_READ_0/chan2_data[5]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[5]\);
    
    HIEFFPLA_INST_0_68203 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\, B => 
        HIEFFPLA_NET_0_72620, C => HIEFFPLA_NET_0_72703, Y => 
        HIEFFPLA_NET_0_72707);
    
    HIEFFPLA_INST_0_55908 : AX1B
      port map(A => HIEFFPLA_NET_0_75418, B => 
        \Communications_0/UART_1/tx_clk_count_i_0[3]\, C => 
        \Communications_0/UART_1/tx_clk_count_i_0[4]\, Y => 
        HIEFFPLA_NET_0_75399);
    
    \Science_0/ADC_READ_0/chan0_data[11]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[17]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[11]\);
    
    HIEFFPLA_INST_0_66833 : NOR3A
      port map(A => HIEFFPLA_NET_0_73021, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73025);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[2]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72337, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[2]_net_1\);
    
    HIEFFPLA_INST_0_61312 : AND2A
      port map(A => HIEFFPLA_NET_0_74217, B => 
        HIEFFPLA_NET_0_74211, Y => HIEFFPLA_NET_0_74220);
    
    \General_Controller_0/st_wdata[11]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[11]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[11]\);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[5]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72334, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[5]_net_1\);
    
    HIEFFPLA_INST_0_70618 : AX1C
      port map(A => HIEFFPLA_NET_0_72070, B => 
        \Timing_0/m_time[4]_net_1\, C => 
        \Timing_0/m_time[5]_net_1\, Y => HIEFFPLA_NET_0_72062);
    
    HIEFFPLA_INST_0_67660 : OA1A
      port map(A => General_Controller_0_en_sensors, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/isSetup_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72831);
    
    HIEFFPLA_INST_0_61337 : AX1
      port map(A => HIEFFPLA_NET_0_74262, B => 
        \General_Controller_0/state_seconds[3]_net_1\, C => 
        \General_Controller_0/state_seconds[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74213);
    
    HIEFFPLA_INST_0_56459 : XNOR3
      port map(A => HIEFFPLA_NET_0_75321, B => 
        HIEFFPLA_NET_0_75318, C => HIEFFPLA_NET_0_75317, Y => 
        HIEFFPLA_NET_0_75276);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_WADDR[6]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75288, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[6]\\\\\);
    
    \Pressure_Signal_Debounce_0/ms_cnt[5]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73489, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[5]_net_1\);
    
    \GS_Readout_0/send[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74716, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74630, Q => 
        \GS_Readout_0_send[1]\);
    
    HIEFFPLA_INST_0_63722 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[7]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_nof_steps[7]_net_1\, S
         => \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73722);
    
    HIEFFPLA_INST_0_58179 : AO1
      port map(A => \Sensors_0_mag_y[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75116, Y => HIEFFPLA_NET_0_74835);
    
    HIEFFPLA_INST_0_55451 : AO1
      port map(A => HIEFFPLA_NET_0_75512, B => 
        \Communications_0/UART_0/tx_count[1]_net_1\, C => 
        HIEFFPLA_NET_0_75508, Y => HIEFFPLA_NET_0_75509);
    
    HIEFFPLA_INST_0_70172 : AOI1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\, 
        B => HIEFFPLA_NET_0_72237, C => HIEFFPLA_NET_0_72269, Y
         => HIEFFPLA_NET_0_72202);
    
    HIEFFPLA_INST_0_65461 : NOR2A
      port map(A => HIEFFPLA_NET_0_73369, B => 
        HIEFFPLA_NET_0_73381, Y => HIEFFPLA_NET_0_73370);
    
    HIEFFPLA_INST_0_60187 : MX2
      port map(A => HIEFFPLA_NET_0_74454, B => 
        HIEFFPLA_NET_0_74533, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74448);
    
    HIEFFPLA_INST_0_57930 : AOI1
      port map(A => \Sensors_0_acc_time[12]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74901, Y => HIEFFPLA_NET_0_74902);
    
    HIEFFPLA_INST_0_69029 : AND2
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0_write_done\, B
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        Y => HIEFFPLA_NET_0_72492);
    
    HIEFFPLA_INST_0_67656 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        B => HIEFFPLA_NET_0_72792, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, Y
         => HIEFFPLA_NET_0_72832);
    
    \Science_0/ADC_READ_0/exp_packet_1[9]\ : DFN1E0
      port map(D => \AFLSDF_INV_11\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[9]\);
    
    HIEFFPLA_INST_0_67253 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        B => HIEFFPLA_NET_0_72761, Y => HIEFFPLA_NET_0_72927);
    
    HIEFFPLA_INST_0_65023 : AO1B
      port map(A => HIEFFPLA_NET_0_73447, B => 
        HIEFFPLA_NET_0_73477, C => HIEFFPLA_NET_0_73482, Y => 
        HIEFFPLA_NET_0_73486);
    
    HIEFFPLA_INST_0_64626 : NAND3C
      port map(A => HIEFFPLA_NET_0_73622, B => 
        HIEFFPLA_NET_0_73555, C => HIEFFPLA_NET_0_73613, Y => 
        HIEFFPLA_NET_0_73582);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/i2c_addr_1[0]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_72480, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72549, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_i2c_addr[0]\);
    
    HIEFFPLA_INST_0_69499 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[2]_net_1\, 
        C => HIEFFPLA_NET_0_72346, Y => HIEFFPLA_NET_0_72376);
    
    HIEFFPLA_INST_0_64682 : NOR3B
      port map(A => HIEFFPLA_NET_0_74039, B => 
        HIEFFPLA_NET_0_73564, C => HIEFFPLA_NET_0_73928, Y => 
        HIEFFPLA_NET_0_73565);
    
    \Timekeeper_0/microseconds[22]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72137, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[22]\);
    
    HIEFFPLA_INST_0_70022 : NAND2
      port map(A => General_Controller_0_en_sensors, B => 
        \Sensors_0/Pressure_Sensor_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72245);
    
    \Science_0/ADC_READ_0/exp_packet_1[70]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[14]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[70]\);
    
    HIEFFPLA_INST_0_68692 : AND3
      port map(A => HIEFFPLA_NET_0_72584, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_we\, C => 
        HIEFFPLA_NET_0_72669, Y => HIEFFPLA_NET_0_72585);
    
    HIEFFPLA_INST_0_69253 : AND2B
      port map(A => \Sensors_0/Gyro_0/state[8]\, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, Y
         => HIEFFPLA_NET_0_72438);
    
    HIEFFPLA_INST_0_62482 : NOR3A
      port map(A => HIEFFPLA_NET_0_73900, B => 
        \General_Controller_0/uc_rx_state_0[1]_net_1\, C => 
        HIEFFPLA_NET_0_73897, Y => HIEFFPLA_NET_0_73973);
    
    HIEFFPLA_INST_0_71012 : AOI1C
      port map(A => \I2C_PassThrough_0/state[0]_net_1\, B => 
        UC_I2C4_SDA_in, C => HIEFFPLA_NET_0_71989, Y => 
        HIEFFPLA_NET_0_73513);
    
    HIEFFPLA_INST_0_57843 : AO1
      port map(A => \Science_0_exp_packet_0[75]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75140, Y => HIEFFPLA_NET_0_74928);
    
    \General_Controller_0/st_waddr[0]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[0]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_waddr[0]\);
    
    CLKINT_1 : CLKINT
      port map(A => RESET_c, Y => CLKINT_1_Y);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[22]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72282, Q => 
        \Sensors_0_pressure_temp_raw[22]\);
    
    HIEFFPLA_INST_0_60588 : MX2
      port map(A => \Science_0_chan7_data[3]\, B => 
        \Science_0_chan7_data[7]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74391);
    
    HIEFFPLA_INST_0_69366 : MX2A
      port map(A => HIEFFPLA_NET_0_72403, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_num_bytes[1]\, 
        S => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72407);
    
    \Science_0/ADC_READ_0/exp_packet_1[58]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[2]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[58]\);
    
    \General_Controller_0/status_bits_1[34]\ : DFN1E1
      port map(D => Eject_Signal_Debounce_0_ffu_ejected_out, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74266, Q => 
        \Data_Hub_Packets_0_status_packet[1]\);
    
    \Science_0/ADC_READ_0/chan4_data[9]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[9]\);
    
    \Pressure_Signal_Debounce_0/ms_cnt[7]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73486, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[7]_net_1\);
    
    \Timekeeper_0/microseconds[13]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72147, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[13]\);
    
    HIEFFPLA_INST_0_67615 : AND3
      port map(A => HIEFFPLA_NET_0_72894, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, C
         => HIEFFPLA_NET_0_72752, Y => HIEFFPLA_NET_0_72842);
    
    HIEFFPLA_INST_0_58246 : AO1
      port map(A => \Sensors_0_gyro_time[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75113, Y => HIEFFPLA_NET_0_74821);
    
    HIEFFPLA_INST_0_61860 : AND3
      port map(A => HIEFFPLA_NET_0_74087, B => 
        HIEFFPLA_NET_0_74107, C => HIEFFPLA_NET_0_73880, Y => 
        HIEFFPLA_NET_0_74114);
    
    HIEFFPLA_INST_0_66861 : AND3
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_we\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73019);
    
    HIEFFPLA_INST_0_55472 : XA1B
      port map(A => \Communications_0/UART_0/tx_state[0]_net_1\, 
        B => \Communications_0/UART_0/tx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_75528, Y => HIEFFPLA_NET_0_75503);
    
    HIEFFPLA_INST_0_67998 : OR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, B
         => HIEFFPLA_NET_0_72744, C => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_72757);
    
    HIEFFPLA_INST_0_70808 : OR3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        Y => HIEFFPLA_NET_0_72008);
    
    HIEFFPLA_INST_0_68738 : NOR3B
      port map(A => HIEFFPLA_NET_0_72701, B => 
        HIEFFPLA_NET_0_72634, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72573);
    
    HIEFFPLA_INST_0_60891 : OR3B
      port map(A => \General_Controller_0/command[1]_net_1\, B
         => \General_Controller_0/command[2]_net_1\, C => 
        \General_Controller_0/command[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74328);
    
    HIEFFPLA_INST_0_66906 : NAND3C
      port map(A => HIEFFPLA_NET_0_72935, B => 
        HIEFFPLA_NET_0_72751, C => HIEFFPLA_NET_0_72762, Y => 
        HIEFFPLA_NET_0_73007);
    
    HIEFFPLA_INST_0_56602 : MX2
      port map(A => HIEFFPLA_NET_0_75200, B => 
        HIEFFPLA_NET_0_75072, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75233);
    
    \Communications_0/UART_1/rx_clk_count[25]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75463, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75443, Q => 
        \Communications_0/UART_1/rx_clk_count[25]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[20]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[20]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[20]\);
    
    \General_Controller_0/sweep_table_nof_steps[5]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73980, Q => 
        \General_Controller_0/sweep_table_nof_steps[5]_net_1\);
    
    \L4WR_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => L4WR_c, E => \VCC\, DOUT => 
        \L4WR_pad/U0/NET1\, EOUT => \L4WR_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_65736 : AND3B
      port map(A => \Science_0/ADC_READ_0/cnt[2]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_73294, Y => HIEFFPLA_NET_0_73295);
    
    HIEFFPLA_INST_0_68587 : AND3C
      port map(A => HIEFFPLA_NET_0_72601, B => 
        HIEFFPLA_NET_0_72596, C => HIEFFPLA_NET_0_72594, Y => 
        HIEFFPLA_NET_0_72611);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[7]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[7]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[7]\);
    
    \Communications_0/UART_0/rx_clk_count[31]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75568, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75554, Q => 
        \Communications_0/UART_0/rx_clk_count_c0\);
    
    HIEFFPLA_INST_0_70373 : AND3
      port map(A => \Timekeeper_0_microseconds[7]\, B => 
        HIEFFPLA_NET_0_72159, C => \Timekeeper_0_microseconds[8]\, 
        Y => HIEFFPLA_NET_0_72157);
    
    HIEFFPLA_INST_0_55843 : AO1
      port map(A => HIEFFPLA_NET_0_75416, B => 
        HIEFFPLA_NET_0_75417, C => 
        \Communications_0/UART_1/tx_clk_count_i_0[4]\, Y => 
        HIEFFPLA_NET_0_75413);
    
    HIEFFPLA_INST_0_68729 : XA1B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\, B
         => \Sensors_0/Gyro_0/I2C_Master_0/next_state[0]_net_1\, 
        C => \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72576);
    
    HIEFFPLA_INST_0_56090 : NOR3B
      port map(A => HIEFFPLA_NET_0_75351, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[7]\\\\\, C
         => HIEFFPLA_NET_0_75373, Y => HIEFFPLA_NET_0_75349);
    
    HIEFFPLA_INST_0_58302 : AO1
      port map(A => \Sensors_0_mag_x[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75106, Y => HIEFFPLA_NET_0_74807);
    
    HIEFFPLA_INST_0_58007 : AO1B
      port map(A => \Sensors_0_mag_time[16]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74880, Y => HIEFFPLA_NET_0_74881);
    
    \General_Controller_0/unit_id[5]\ : DFN1E0P1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, PRE => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73990, Q => 
        \General_Controller_0_unit_id[5]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[50]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[16]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[50]\);
    
    \I2C_PassThrough_0/cnt[2]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73517, CLK => CLKINT_0_Y_0, Q
         => \I2C_PassThrough_0/cnt[2]_net_1\);
    
    HIEFFPLA_INST_0_68022 : NAND3C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72752);
    
    HIEFFPLA_INST_0_58607 : AND2B
      port map(A => \GS_Readout_0/prevState[4]_net_1\, B => 
        \GS_Readout_0/prevState[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74721);
    
    \General_Controller_0/sweep_table_sweep_cnt[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74134, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[4]_net_1\);
    
    HIEFFPLA_INST_0_69382 : AND3A
      port map(A => HIEFFPLA_NET_0_72426, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        C => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72402);
    
    HIEFFPLA_INST_0_70883 : AX1E
      port map(A => HIEFFPLA_NET_0_72711, B => 
        HIEFFPLA_NET_0_72876, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72005);
    
    HIEFFPLA_INST_0_56215 : OR2A
      port map(A => \Data_Saving_0/Packet_Saver_0_we\, B => 
        \Data_Saving_0/FPGA_Buffer_0/full\, Y => 
        \Data_Saving_0/FPGA_Buffer_0/MEMWENEG\);
    
    HIEFFPLA_INST_0_61891 : MX2A
      port map(A => \General_Controller_0/uc_rx_byte[3]_net_1\, B
         => \General_Controller_0/uc_rx_byte[0]_net_1\, S => 
        \General_Controller_0/uc_rx_byte[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74108);
    
    HIEFFPLA_INST_0_65768 : AND2A
      port map(A => HIEFFPLA_NET_0_73241, B => 
        HIEFFPLA_NET_0_73283, Y => HIEFFPLA_NET_0_73284);
    
    HIEFFPLA_INST_0_58499 : NAND3C
      port map(A => HIEFFPLA_NET_0_74750, B => 
        \Eject_Signal_Debounce_0/ms_cnt[2]_net_1\, C => 
        \Eject_Signal_Debounce_0/ms_cnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74748);
    
    HIEFFPLA_INST_0_56504 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, B
         => HIEFFPLA_NET_0_75352, Y => HIEFFPLA_NET_0_75261);
    
    \FMC_DA_pad[1]/U0/U1\ : IOTRI_OB_EB
      port map(D => \FMC_DA_c[1]\, E => \VCC\, DOUT => 
        \FMC_DA_pad[1]/U0/NET1\, EOUT => \FMC_DA_pad[1]/U0/NET2\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[9]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[9]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[9]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[6]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72482, Q => 
        \Sensors_0_gyro_y[6]\);
    
    HIEFFPLA_INST_0_66059 : NAND2
      port map(A => \Science_0/DAC_SET_0/cnt[1]_net_1\, B => 
        \Science_0/DAC_SET_0/cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73223);
    
    HIEFFPLA_INST_0_66742 : AND3
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        B => ACCE_SDA_in, C => ACCE_SCL_c, Y => 
        HIEFFPLA_NET_0_73048);
    
    \Science_0/ADC_READ_0/cnt4up[2]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73304, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4up[2]_net_1\);
    
    HIEFFPLA_INST_0_68259 : XAI1A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, B => 
        HIEFFPLA_NET_0_72572, C => HIEFFPLA_NET_0_72622, Y => 
        HIEFFPLA_NET_0_72695);
    
    AFLSDF_INV_34 : INV
      port map(A => CLKINT_1_Y, Y => \AFLSDF_INV_34\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/temp[1]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72555, Q => 
        \Sensors_0_gyro_temp[1]\);
    
    HIEFFPLA_INST_0_70309 : NOR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        Y => HIEFFPLA_NET_0_72177);
    
    HIEFFPLA_INST_0_59569 : MX2
      port map(A => HIEFFPLA_NET_0_74476, B => 
        HIEFFPLA_NET_0_74366, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74536);
    
    HIEFFPLA_INST_0_60097 : MX2
      port map(A => HIEFFPLA_NET_0_74471, B => 
        HIEFFPLA_NET_0_74530, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74462);
    
    HIEFFPLA_INST_0_56520 : AND3
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[5]_net_1\, B
         => HIEFFPLA_NET_0_75254, C => 
        \Data_Saving_0/Interrupt_Generator_0/counter[6]_net_1\, Y
         => HIEFFPLA_NET_0_75255);
    
    HIEFFPLA_INST_0_57605 : AO1B
      port map(A => \Sensors_0_gyro_x[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74994, Y => HIEFFPLA_NET_0_74995);
    
    \Science_0/ADC_READ_0/chan5_data[2]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[2]\);
    
    HIEFFPLA_INST_0_70692 : AX1C
      port map(A => HIEFFPLA_NET_0_72039, B => 
        \Timing_0/s_time[6]_net_1\, C => 
        \Timing_0/s_time[7]_net_1\, Y => HIEFFPLA_NET_0_72042);
    
    HIEFFPLA_INST_0_60956 : NAND3C
      port map(A => HIEFFPLA_NET_0_74310, B => 
        \Timekeeper_0_milliseconds[9]\, C => 
        \Timekeeper_0_milliseconds[7]\, Y => HIEFFPLA_NET_0_74311);
    
    \General_Controller_0/sweep_table_write_value[15]\ : DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[15]_net_1\);
    
    HIEFFPLA_INST_0_57657 : AO1
      port map(A => \Sensors_0_pressure_raw[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74792, Y => HIEFFPLA_NET_0_74979);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRYSYNC[8]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_17_Q\, 
        CLK => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[8]\\\\\);
    
    HIEFFPLA_INST_0_54954 : AX1C
      port map(A => \ClockDivs_0/cnt_800kHz[0]_net_1\, B => 
        \ClockDivs_0/cnt_800kHz[1]_net_1\, C => 
        \ClockDivs_0/cnt_800kHz[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75629);
    
    HIEFFPLA_INST_0_56236 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[8]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[7]\\\\\, Y => 
        HIEFFPLA_NET_0_75328);
    
    \General_Controller_0/sweep_table_probe_id[2]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73924, Q => 
        \General_Controller_0/sweep_table_probe_id[2]_net_1\);
    
    \Science_0/ADC_READ_0/data_a[0]\ : DFN1E1C1
      port map(D => AB_c, CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, 
        E => \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[0]_net_1\);
    
    HIEFFPLA_INST_0_66435 : AND3A
      port map(A => HIEFFPLA_NET_0_73121, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73122);
    
    HIEFFPLA_INST_0_70353 : AND3
      port map(A => \Timekeeper_0_microseconds[15]\, B => 
        HIEFFPLA_NET_0_72161, C => 
        \Timekeeper_0_microseconds[16]\, Y => 
        HIEFFPLA_NET_0_72162);
    
    HIEFFPLA_INST_0_67423 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, 
        Y => HIEFFPLA_NET_0_72885);
    
    HIEFFPLA_INST_0_61681 : MX2
      port map(A => \SweepTable_0_RD[3]\, B => 
        \SweepTable_1_RD[3]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74161);
    
    HIEFFPLA_INST_0_55706 : AOI1B
      port map(A => HIEFFPLA_NET_0_75481, B => 
        HIEFFPLA_NET_0_75479, C => HIEFFPLA_NET_0_75440, Y => 
        HIEFFPLA_NET_0_75441);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[0]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[0]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[0]\);
    
    HIEFFPLA_INST_0_59421 : MX2
      port map(A => HIEFFPLA_NET_0_74506, B => 
        HIEFFPLA_NET_0_74357, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74556);
    
    HIEFFPLA_INST_0_56291 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[4]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[3]\\\\\, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[2]\\\\\, Y => 
        HIEFFPLA_NET_0_75317);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72467, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[2]_net_1\);
    
    HIEFFPLA_INST_0_69355 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72409);
    
    HIEFFPLA_INST_0_61794 : XOR2
      port map(A => HIEFFPLA_NET_0_74146, B => 
        \General_Controller_0/sweep_table_sweep_cnt[9]_net_1\, Y
         => HIEFFPLA_NET_0_74129);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[4]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72800, Q => 
        \Sensors_0_acc_x[4]\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[2]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75265, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[2]\\\\\);
    
    HIEFFPLA_INST_0_61570 : AND3C
      port map(A => 
        \General_Controller_0/sweep_table_probe_id[3]_net_1\, B
         => \General_Controller_0/sweep_table_probe_id[2]_net_1\, 
        C => \General_Controller_0/sweep_table_probe_id[1]_net_1\, 
        Y => HIEFFPLA_NET_0_74182);
    
    HIEFFPLA_INST_0_64458 : OA1C
      port map(A => HIEFFPLA_NET_0_73592, B => 
        \General_Controller_0/uc_tx_state[0]_net_1\, C => 
        HIEFFPLA_NET_0_73560, Y => HIEFFPLA_NET_0_73622);
    
    HIEFFPLA_INST_0_64730 : MX2A
      port map(A => Communications_0_uc_tx_rdy, B => 
        HIEFFPLA_NET_0_73529, S => HIEFFPLA_NET_0_73521, Y => 
        HIEFFPLA_NET_0_73551);
    
    HIEFFPLA_INST_0_68220 : AND3C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72702);
    
    HIEFFPLA_INST_0_64169 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_1[7]_net_1\, 
        B => 
        \General_Controller_0/constant_bias_voltage_1[15]_net_1\, 
        S => \General_Controller_0/uc_tx_substate[1]_net_1\, Y
         => HIEFFPLA_NET_0_73658);
    
    \Data_Saving_0/Packet_Saver_0/data_out[8]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75205, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[8]\);
    
    \Communications_0/UART_1/rx_rdy\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75444, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75446, Q => 
        Communications_0_uc_rx_rdy);
    
    HIEFFPLA_INST_0_64653 : AND2
      port map(A => 
        \General_Controller_0/uc_tx_nextstate[0]_net_1\, B => 
        HIEFFPLA_NET_0_73584, Y => HIEFFPLA_NET_0_73575);
    
    \Science_0/ADC_READ_0/chan6_data[3]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[3]\);
    
    \Science_0/ADC_READ_0/chan0_data[3]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[3]\);
    
    HIEFFPLA_INST_0_69526 : AOI1D
      port map(A => HIEFFPLA_NET_0_72366, B => 
        HIEFFPLA_NET_0_72365, C => HIEFFPLA_NET_0_72350, Y => 
        HIEFFPLA_NET_0_72371);
    
    HIEFFPLA_INST_0_57512 : AOI1
      port map(A => \Science_0_exp_packet_0[21]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_75023, Y => HIEFFPLA_NET_0_75024);
    
    HIEFFPLA_INST_0_70071 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]_net_1\, 
        B => HIEFFPLA_NET_0_72237, C => HIEFFPLA_NET_0_72222, Y
         => HIEFFPLA_NET_0_72229);
    
    HIEFFPLA_INST_0_58010 : AOI1
      port map(A => \Sensors_0_acc_time[16]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74879, Y => HIEFFPLA_NET_0_74880);
    
    HIEFFPLA_INST_0_66382 : OR3A
      port map(A => HIEFFPLA_NET_0_73042, B => 
        HIEFFPLA_NET_0_73059, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73133);
    
    HIEFFPLA_INST_0_68217 : NAND3
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72703);
    
    HIEFFPLA_INST_0_70151 : AND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72208);
    
    \General_Controller_0/sweep_table_points[4]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[4]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[4]_net_1\);
    
    \General_Controller_0/sweep_table_points[0]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[0]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[0]_net_1\);
    
    HIEFFPLA_INST_0_67354 : OR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72900);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[13]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72484, Q => 
        \Sensors_0_gyro_y[13]\);
    
    \Science_0/DAC_SET_0/cnt[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73216, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/cnt[3]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/i2c_addr_1[2]\ : 
        DFN1E0
      port map(D => HIEFFPLA_NET_0_72991, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72774, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[2]\);
    
    HIEFFPLA_INST_0_63260 : NOR3B
      port map(A => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, B => 
        HIEFFPLA_NET_0_73905, C => HIEFFPLA_NET_0_73869, Y => 
        HIEFFPLA_NET_0_73797);
    
    HIEFFPLA_INST_0_69013 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        B => HIEFFPLA_NET_0_72540, C => HIEFFPLA_NET_0_72497, Y
         => HIEFFPLA_NET_0_72498);
    
    HIEFFPLA_INST_0_62531 : OR3A
      port map(A => HIEFFPLA_NET_0_74091, B => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, C => 
        HIEFFPLA_NET_0_74119, Y => HIEFFPLA_NET_0_73963);
    
    HIEFFPLA_INST_0_68377 : AO1
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, C => 
        HIEFFPLA_NET_0_72630, Y => HIEFFPLA_NET_0_72665);
    
    \Science_0/ADC_READ_0/data_b[2]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[1]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[2]_net_1\);
    
    \General_Controller_0/sweep_table_sweep_cnt[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74137, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[1]_net_1\);
    
    \General_Controller_0/sweep_table_step_id[6]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73926, Q => 
        \General_Controller_0/sweep_table_step_id[6]_net_1\);
    
    \LDCLK_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => LDCLK_c, E => \VCC\, DOUT => 
        \LDCLK_pad/U0/NET1\, EOUT => \LDCLK_pad/U0/NET2\);
    
    \FMC_DA_pad[5]/U0/U0\ : IOPAD_TRI
      port map(D => \FMC_DA_pad[5]/U0/NET1\, E => 
        \FMC_DA_pad[5]/U0/NET2\, PAD => FMC_DA(5));
    
    \General_Controller_0/state_seconds[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74222, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[5]_net_1\);
    
    HIEFFPLA_INST_0_70332 : AND2
      port map(A => HIEFFPLA_NET_0_72232, B => 
        \Sensors_0/Pressure_Sensor_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72172);
    
    HIEFFPLA_INST_0_55120 : AND2B
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[29]_net_1\, B => 
        \Communications_0/UART_0/rx_clk_count[30]_net_1\, Y => 
        HIEFFPLA_NET_0_75584);
    
    HIEFFPLA_INST_0_63277 : AND3
      port map(A => HIEFFPLA_NET_0_73900, B => 
        HIEFFPLA_NET_0_73906, C => HIEFFPLA_NET_0_73796, Y => 
        HIEFFPLA_NET_0_73792);
    
    HIEFFPLA_INST_0_59181 : NOR3A
      port map(A => \GS_Readout_0/state[0]_net_1\, B => 
        Communications_0_ext_tx_rdy, C => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74594);
    
    HIEFFPLA_INST_0_55565 : AO1C
      port map(A => \Communications_0/UART_1/rx_clk_count_c0\, B
         => HIEFFPLA_NET_0_75471, C => 
        \Communications_0/UART_1/rx_clk_count[28]_net_1\, Y => 
        HIEFFPLA_NET_0_75479);
    
    HIEFFPLA_INST_0_67098 : AO1A
      port map(A => HIEFFPLA_NET_0_72761, B => 
        HIEFFPLA_NET_0_72934, C => HIEFFPLA_NET_0_72766, Y => 
        HIEFFPLA_NET_0_72964);
    
    HIEFFPLA_INST_0_65379 : XOR2
      port map(A => \Science_0/ADC_READ_0/cnt1up[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt1up[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73395);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_19\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[8]\\\\\, CLK => 
        CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_19_Q\);
    
    HIEFFPLA_INST_0_62427 : AND3
      port map(A => HIEFFPLA_NET_0_73777, B => 
        HIEFFPLA_NET_0_74171, C => HIEFFPLA_NET_0_73972, Y => 
        HIEFFPLA_NET_0_73984);
    
    HIEFFPLA_INST_0_62246 : NOR3A
      port map(A => HIEFFPLA_NET_0_73991, B => 
        HIEFFPLA_NET_0_73804, C => HIEFFPLA_NET_0_73788, Y => 
        HIEFFPLA_NET_0_74021);
    
    HIEFFPLA_INST_0_65689 : AO1A
      port map(A => HIEFFPLA_NET_0_73308, B => 
        HIEFFPLA_NET_0_73276, C => HIEFFPLA_NET_0_73422, Y => 
        HIEFFPLA_NET_0_73309);
    
    \General_Controller_0/status_bits_1[55]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74191, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[55]\);
    
    AFLSDF_INV_19 : INV
      port map(A => \m_time[7]\, Y => \AFLSDF_INV_19\);
    
    HIEFFPLA_INST_0_67700 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, 
        Y => HIEFFPLA_NET_0_72820);
    
    HIEFFPLA_INST_0_59775 : NOR2A
      port map(A => HIEFFPLA_NET_0_74439, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74510);
    
    HIEFFPLA_INST_0_62303 : NOR2A
      port map(A => \General_Controller_0/uc_rx_state[3]_net_1\, 
        B => HIEFFPLA_NET_0_73781, Y => HIEFFPLA_NET_0_74010);
    
    HIEFFPLA_INST_0_66503 : AND2
      port map(A => HIEFFPLA_NET_0_73132, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73107);
    
    \Science_0/ADC_READ_0/exp_packet_1[27]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[11]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[27]\);
    
    HIEFFPLA_INST_0_70033 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[2]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72240);
    
    \ACCE_SCL_pad/U0/U0\ : IOPAD_TRI
      port map(D => \ACCE_SCL_pad/U0/NET1\, E => 
        \ACCE_SCL_pad/U0/NET2\, PAD => ACCE_SCL);
    
    HIEFFPLA_INST_0_64739 : MX2
      port map(A => HIEFFPLA_NET_0_73548, B => 
        HIEFFPLA_NET_0_73531, S => HIEFFPLA_NET_0_73521, Y => 
        HIEFFPLA_NET_0_73550);
    
    HIEFFPLA_INST_0_61058 : AO1C
      port map(A => Eject_Signal_Debounce_0_ffu_ejected_out, B
         => \General_Controller_0/flight_state[2]_net_1\, C => 
        HIEFFPLA_NET_0_74296, Y => HIEFFPLA_NET_0_74285);
    
    HIEFFPLA_INST_0_68715 : AO1A
      port map(A => HIEFFPLA_NET_0_72577, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, C
         => HIEFFPLA_NET_0_72579, Y => HIEFFPLA_NET_0_72580);
    
    HIEFFPLA_INST_0_66701 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73059);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[0]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[0]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[0]\);
    
    HIEFFPLA_INST_0_68077 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72736);
    
    HIEFFPLA_INST_0_67128 : AND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72959);
    
    AFLSDF_INV_17 : INV
      port map(A => HIEFFPLA_NET_0_72494, Y => \AFLSDF_INV_17\);
    
    \Timekeeper_0/microseconds[10]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72150, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[10]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[21]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[21]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[21]\);
    
    \GS_Readout_0/send[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74713, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74630, Q => 
        \GS_Readout_0_send[4]\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[10]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75267, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[10]\\\\\);
    
    HIEFFPLA_INST_0_55298 : MX2
      port map(A => HIEFFPLA_NET_0_75542, B => 
        HIEFFPLA_NET_0_75541, S => 
        \Communications_0/UART_0/tx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75543);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/scl\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_72379, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        PRESSURE_SCL_c);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[6]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72804, Q => 
        \Sensors_0_mag_x[6]\);
    
    HIEFFPLA_INST_0_64803 : AND2
      port map(A => 
        \General_Controller_0/sweep_table_write_wait[0]_net_1\, B
         => HIEFFPLA_NET_0_74127, Y => HIEFFPLA_NET_0_73538);
    
    \Science_0/DAC_SET_0/state[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73210, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/state[3]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[72]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[16]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[72]\);
    
    HIEFFPLA_INST_0_69408 : AND3
      port map(A => HIEFFPLA_NET_0_72351, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        C => HIEFFPLA_NET_0_72428, Y => HIEFFPLA_NET_0_72396);
    
    HIEFFPLA_INST_0_69829 : XA1A
      port map(A => HIEFFPLA_NET_0_72309, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[6]_net_1\, 
        C => HIEFFPLA_NET_0_72236, Y => HIEFFPLA_NET_0_72293);
    
    HIEFFPLA_INST_0_70974 : MX2A
      port map(A => HIEFFPLA_NET_0_71996, B => 
        \Science_0/ADC_READ_0_G4[1]\, S => HIEFFPLA_NET_0_73319, 
        Y => HIEFFPLA_NET_0_73249);
    
    HIEFFPLA_INST_0_56023 : AND3
      port map(A => HIEFFPLA_NET_0_75375, B => 
        HIEFFPLA_NET_0_75364, C => HIEFFPLA_NET_0_75366, Y => 
        HIEFFPLA_NET_0_75367);
    
    \Timekeeper_0/milliseconds[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72098, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[4]\);
    
    \General_Controller_0/sweep_table_samples_per_point[2]\ : 
        DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[2]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[2]_net_1\);
    
    HIEFFPLA_INST_0_68264 : XA1
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\, B => 
        HIEFFPLA_NET_0_72573, C => HIEFFPLA_NET_0_72622, Y => 
        HIEFFPLA_NET_0_72694);
    
    \Timekeeper_0/milliseconds[17]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72108, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[17]\);
    
    HIEFFPLA_INST_0_61342 : NOR2A
      port map(A => \General_Controller_0/state_seconds[5]_net_1\, 
        B => HIEFFPLA_NET_0_74248, Y => HIEFFPLA_NET_0_74212);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[15]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[15]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[15]\);
    
    HIEFFPLA_INST_0_69371 : XA1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[2]_net_1\, 
        B => HIEFFPLA_NET_0_72409, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72406);
    
    HIEFFPLA_INST_0_56517 : AND3
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[1]_net_1\, B
         => 
        \Data_Saving_0/Interrupt_Generator_0/counter[0]_net_1\, C
         => 
        \Data_Saving_0/Interrupt_Generator_0/counter[2]_net_1\, Y
         => HIEFFPLA_NET_0_75256);
    
    HIEFFPLA_INST_0_55973 : AO1
      port map(A => TOP_UART_RX_c, B => EMU_RX_c, C => 
        UC_CONSOLE_EN_c, Y => HIEFFPLA_NET_0_75380);
    
    HIEFFPLA_INST_0_65997 : AND2B
      port map(A => \Science_0/ADC_READ_0_G4[0]\, B => 
        \Science_0/ADC_READ_0_G4[1]\, Y => HIEFFPLA_NET_0_73245);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[8]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72782, Q => 
        \Sensors_0_mag_y[8]\);
    
    HIEFFPLA_INST_0_88373 : XA1B
      port map(A => HIEFFPLA_NET_0_75288, B => 
        HIEFFPLA_NET_0_75321, C => HIEFFPLA_NET_0_88383, Y => 
        HIEFFPLA_NET_0_88386);
    
    HIEFFPLA_INST_0_69386 : NOR3A
      port map(A => HIEFFPLA_NET_0_72351, B => 
        HIEFFPLA_NET_0_72423, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72401);
    
    \General_Controller_0/st_ren0\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74176, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74174, Q => 
        \SweepTable_0/WEBP\);
    
    HIEFFPLA_INST_0_62912 : NAND3C
      port map(A => HIEFFPLA_NET_0_73877, B => 
        HIEFFPLA_NET_0_73813, C => HIEFFPLA_NET_0_74043, Y => 
        HIEFFPLA_NET_0_73867);
    
    HIEFFPLA_INST_0_70535 : AND3
      port map(A => \Timing_0/f_time[0]_net_1\, B => 
        \Timing_0/f_time[1]_net_1\, C => 
        \Timing_0/f_time[2]_net_1\, Y => HIEFFPLA_NET_0_72090);
    
    HIEFFPLA_INST_0_58885 : AOI1
      port map(A => HIEFFPLA_NET_0_74693, B => 
        HIEFFPLA_NET_0_74499, C => HIEFFPLA_NET_0_74665, Y => 
        HIEFFPLA_NET_0_74666);
    
    HIEFFPLA_INST_0_65801 : AO16
      port map(A => \Science_0/ADC_READ_0/data_b[15]_net_1\, B
         => \Science_0/ADC_READ_0/data_b[16]_net_1\, C => 
        \Science_0/ADC_READ_0/data_b[17]_net_1\, Y => 
        HIEFFPLA_NET_0_73277);
    
    HIEFFPLA_INST_0_55729 : MX2
      port map(A => HIEFFPLA_NET_0_75434, B => 
        HIEFFPLA_NET_0_75432, S => 
        \Communications_0/UART_1/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75436);
    
    \General_Controller_0/sweep_table_points[11]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[11]_net_1\);
    
    HIEFFPLA_INST_0_68763 : NAND3C
      port map(A => HIEFFPLA_NET_0_72565, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, C
         => HIEFFPLA_NET_0_72550, Y => HIEFFPLA_NET_0_72567);
    
    HIEFFPLA_INST_0_67002 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[3]\, 
        C => HIEFFPLA_NET_0_72884, Y => HIEFFPLA_NET_0_72987);
    
    HIEFFPLA_INST_0_58921 : AND3C
      port map(A => HIEFFPLA_NET_0_74624, B => 
        HIEFFPLA_NET_0_74657, C => HIEFFPLA_NET_0_74618, Y => 
        HIEFFPLA_NET_0_74658);
    
    \General_Controller_0/uc_tx_state[14]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73938, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[14]_net_1\);
    
    HIEFFPLA_INST_0_68083 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72734);
    
    HIEFFPLA_INST_0_57608 : AOI1
      port map(A => \Science_0_exp_packet_0[45]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74800, Y => HIEFFPLA_NET_0_74994);
    
    HIEFFPLA_INST_0_66478 : AOI1D
      port map(A => HIEFFPLA_NET_0_73109, B => 
        HIEFFPLA_NET_0_73112, C => HIEFFPLA_NET_0_73065, Y => 
        HIEFFPLA_NET_0_73110);
    
    HIEFFPLA_INST_0_70114 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        B => HIEFFPLA_NET_0_72269, C => HIEFFPLA_NET_0_72208, Y
         => HIEFFPLA_NET_0_72215);
    
    HIEFFPLA_INST_0_61149 : AND3C
      port map(A => \General_Controller_0/state_seconds[0]_net_1\, 
        B => \General_Controller_0/state_seconds[2]_net_1\, C => 
        \General_Controller_0/state_seconds[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74263);
    
    HIEFFPLA_INST_0_55110 : NAND3C
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[24]_net_1\, B => 
        \Communications_0/UART_0/rx_clk_count[25]_net_1\, C => 
        \Communications_0/UART_0/rx_clk_count[26]_net_1\, Y => 
        HIEFFPLA_NET_0_75587);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[19]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[19]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[19]\);
    
    HIEFFPLA_INST_0_62355 : NAND3C
      port map(A => HIEFFPLA_NET_0_73929, B => 
        HIEFFPLA_NET_0_73806, C => HIEFFPLA_NET_0_73980, Y => 
        HIEFFPLA_NET_0_73998);
    
    HIEFFPLA_INST_0_69691 : AO1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_we\, 
        C => HIEFFPLA_NET_0_72324, Y => HIEFFPLA_NET_0_72328);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_afull\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75347, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0_afull\);
    
    \Science_0/ADC_READ_0/chan7_data[3]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[3]\);
    
    HIEFFPLA_INST_0_55358 : AO1
      port map(A => HIEFFPLA_NET_0_75532, B => 
        HIEFFPLA_NET_0_75533, C => 
        \Communications_0/UART_0/tx_clk_count_i_0[4]\, Y => 
        HIEFFPLA_NET_0_75530);
    
    HIEFFPLA_INST_0_65627 : NOR3A
      port map(A => HIEFFPLA_NET_0_73323, B => 
        \Science_0/ADC_READ_0/cnt4dn[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt4dn[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73325);
    
    \General_Controller_0/flight_state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74292, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/flight_state[0]_net_1\);
    
    HIEFFPLA_INST_0_65397 : AND2
      port map(A => HIEFFPLA_NET_0_73388, B => 
        \Science_0/ADC_READ_0/cnt1up[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73389);
    
    HIEFFPLA_INST_0_65307 : AND3
      port map(A => HIEFFPLA_NET_0_73417, B => 
        HIEFFPLA_NET_0_73412, C => HIEFFPLA_NET_0_73277, Y => 
        HIEFFPLA_NET_0_73415);
    
    \Science_0/ADC_READ_0/exp_packet_1[52]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73272, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[52]\);
    
    HIEFFPLA_INST_0_58863 : OR3B
      port map(A => HIEFFPLA_NET_0_74410, B => 
        \GS_Readout_0/state[3]_net_1\, C => HIEFFPLA_NET_0_74725, 
        Y => HIEFFPLA_NET_0_74671);
    
    \General_Controller_0/sweep_table_write_value[8]\ : DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[0]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[8]_net_1\);
    
    HIEFFPLA_INST_0_70954 : NAND3C
      port map(A => HIEFFPLA_NET_0_72001, B => 
        HIEFFPLA_NET_0_72995, C => HIEFFPLA_NET_0_72002, Y => 
        HIEFFPLA_NET_0_72996);
    
    HIEFFPLA_INST_0_70608 : AX1C
      port map(A => HIEFFPLA_NET_0_72069, B => \s_clks_net_0[9]\, 
        C => \Timing_0/m_time[3]_net_1\, Y => 
        HIEFFPLA_NET_0_72066);
    
    HIEFFPLA_INST_0_55113 : NOR3B
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[28]_net_1\, B => 
        \Communications_0/UART_0/rx_clk_count[27]_net_1\, C => 
        HIEFFPLA_NET_0_75579, Y => HIEFFPLA_NET_0_75586);
    
    HIEFFPLA_INST_0_65794 : AO1A
      port map(A => \Science_0/ADC_READ_0/countere\, B => 
        HIEFFPLA_NET_0_73236, C => HIEFFPLA_NET_0_73280, Y => 
        HIEFFPLA_NET_0_73278);
    
    \LA0_pad/U0/U0\ : IOPAD_TRI
      port map(D => \LA0_pad/U0/NET1\, E => \LA0_pad/U0/NET2\, 
        PAD => LA0);
    
    HIEFFPLA_INST_0_65704 : AND2
      port map(A => HIEFFPLA_NET_0_73309, B => 
        HIEFFPLA_NET_0_73303, Y => HIEFFPLA_NET_0_73304);
    
    HIEFFPLA_INST_0_66204 : XOR2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G1[0]_net_1\, B
         => \Science_0/ADC_READ_0_G1[0]\, Y => 
        HIEFFPLA_NET_0_73178);
    
    HIEFFPLA_INST_0_62778 : AND3C
      port map(A => \General_Controller_0/uc_rx_state[1]_net_1\, 
        B => \General_Controller_0/uc_rx_substate[4]_net_1\, C
         => \General_Controller_0/uc_rx_substate[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73907);
    
    \General_Controller_0/status_bits_1[56]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74190, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[56]\);
    
    \Communications_0/UART_1/rx_byte[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75378, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75489, Q => 
        \Communications_0/UART_1/rx_byte[7]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[23]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72280, Q => \Sensors_0_pressure_raw[23]\);
    
    \General_Controller_0/sweep_table_sample_skip[10]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[10]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRYSYNC[2]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_9_Q\, CLK
         => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[2]\\\\\);
    
    HIEFFPLA_INST_0_66592 : MX2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[0]\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[4]\, 
        S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73087);
    
    HIEFFPLA_INST_0_66386 : NAND2B
      port map(A => HIEFFPLA_NET_0_73131, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[3]_net_1\, 
        Y => HIEFFPLA_NET_0_73132);
    
    HIEFFPLA_INST_0_57611 : AO1
      port map(A => \Sensors_0_pressure_raw[14]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74992, Y => HIEFFPLA_NET_0_74993);
    
    \Timekeeper_0/milliseconds[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72097, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[5]\);
    
    HIEFFPLA_INST_0_59357 : MX2
      port map(A => HIEFFPLA_NET_0_74571, B => 
        HIEFFPLA_NET_0_74528, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74564);
    
    HIEFFPLA_INST_0_61750 : AND3
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[11]_net_1\, B
         => HIEFFPLA_NET_0_74149, C => 
        \General_Controller_0/sweep_table_sweep_cnt[12]_net_1\, Y
         => HIEFFPLA_NET_0_74147);
    
    HIEFFPLA_INST_0_60773 : MX2
      port map(A => \ch3_data_net_0[0]\, B => \ch3_data_net_0[4]\, 
        S => \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74361);
    
    \Science_0/ADC_READ_0/chan2_data[10]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[10]\);
    
    HIEFFPLA_INST_0_63668 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[14]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_samples_per_point[14]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73731);
    
    HIEFFPLA_INST_0_58777 : NAND3C
      port map(A => HIEFFPLA_NET_0_74686, B => 
        HIEFFPLA_NET_0_74680, C => HIEFFPLA_NET_0_74663, Y => 
        HIEFFPLA_NET_0_74687);
    
    \General_Controller_0/state_seconds[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74225, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[3]_net_1\);
    
    HIEFFPLA_INST_0_67200 : OR3B
      port map(A => HIEFFPLA_NET_0_72953, B => 
        HIEFFPLA_NET_0_72954, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72941);
    
    \L4WR_pad/U0/U0\ : IOPAD_TRI
      port map(D => \L4WR_pad/U0/NET1\, E => \L4WR_pad/U0/NET2\, 
        PAD => L4WR);
    
    HIEFFPLA_INST_0_64822 : XOR2
      port map(A => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, B => 
        HIEFFPLA_NET_0_73532, Y => HIEFFPLA_NET_0_73531);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[2]\ : 
        DFN0E1
      port map(D => HIEFFPLA_NET_0_72386, CLK => 
        ClockDivs_0_clk_800kHz, E => HIEFFPLA_NET_0_72354, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[2]_net_1\);
    
    HIEFFPLA_INST_0_60805 : NAND3C
      port map(A => HIEFFPLA_NET_0_74548, B => 
        HIEFFPLA_NET_0_74355, C => HIEFFPLA_NET_0_74349, Y => 
        HIEFFPLA_NET_0_74356);
    
    HIEFFPLA_INST_0_67246 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72929);
    
    HIEFFPLA_INST_0_63282 : AND3
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[1]_net_1\, C => 
        HIEFFPLA_NET_0_73789, Y => HIEFFPLA_NET_0_73790);
    
    HIEFFPLA_INST_0_69642 : AO1A
      port map(A => PRESSURE_SCL_c, B => HIEFFPLA_NET_0_72331, C
         => HIEFFPLA_NET_0_72326, Y => HIEFFPLA_NET_0_72338);
    
    HIEFFPLA_INST_0_68131 : MX2
      port map(A => HIEFFPLA_NET_0_72722, B => 
        HIEFFPLA_NET_0_72712, S => HIEFFPLA_NET_0_72876, Y => 
        HIEFFPLA_NET_0_72726);
    
    HIEFFPLA_INST_0_55413 : XO1A
      port map(A => HIEFFPLA_NET_0_75535, B => 
        \Communications_0/UART_0/tx_clk_count_i_0[7]\, C => 
        HIEFFPLA_NET_0_75527, Y => HIEFFPLA_NET_0_75519);
    
    HIEFFPLA_INST_0_61176 : NAND3C
      port map(A => HIEFFPLA_NET_0_74264, B => 
        \General_Controller_0/state_seconds[13]_net_1\, C => 
        HIEFFPLA_NET_0_74256, Y => HIEFFPLA_NET_0_74258);
    
    \Pressure_Signal_Debounce_0/low_pressure\ : DFN1C1
      port map(D => \Pressure_Signal_Debounce_0/state[1]_net_1\, 
        CLK => \m_time[7]\, CLR => CLKINT_1_Y, Q => 
        Pressure_Signal_Debounce_0_low_pressure);
    
    HIEFFPLA_INST_0_70778 : OR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[6]_net_1\, 
        B => HIEFFPLA_NET_0_72309, Y => HIEFFPLA_NET_0_72014);
    
    HIEFFPLA_INST_0_70223 : AO1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[3]_net_1\, 
        B => HIEFFPLA_NET_0_72278, C => HIEFFPLA_NET_0_72312, Y
         => HIEFFPLA_NET_0_72192);
    
    \Communications_0/UART_0/tx_clk_count[3]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75523, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_clk_count_i_0[3]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[35]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[1]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[35]\);
    
    HIEFFPLA_INST_0_71213 : AOI1A
      port map(A => \Communications_0/UART_0/rx_state[1]_net_1\, 
        B => HIEFFPLA_NET_0_75555, C => HIEFFPLA_NET_0_71972, Y
         => HIEFFPLA_NET_0_75561);
    
    HIEFFPLA_INST_0_65505 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt2up[3]_net_1\, B => 
        HIEFFPLA_NET_0_73367, C => HIEFFPLA_NET_0_73366, Y => 
        HIEFFPLA_NET_0_73360);
    
    HIEFFPLA_INST_0_69662 : NAND3C
      port map(A => HIEFFPLA_NET_0_72329, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        C => HIEFFPLA_NET_0_72348, Y => HIEFFPLA_NET_0_72334);
    
    HIEFFPLA_INST_0_67471 : AO1A
      port map(A => HIEFFPLA_NET_0_72855, B => 
        HIEFFPLA_NET_0_72743, C => HIEFFPLA_NET_0_72869, Y => 
        HIEFFPLA_NET_0_72870);
    
    HIEFFPLA_INST_0_65340 : XA1B
      port map(A => HIEFFPLA_NET_0_73410, B => 
        \Science_0/ADC_READ_0/cnt1dn[3]_net_1\, C => 
        HIEFFPLA_NET_0_73244, Y => HIEFFPLA_NET_0_73405);
    
    HIEFFPLA_INST_0_58870 : AND2
      port map(A => \General_Controller_0_gs_id[1]\, B => 
        HIEFFPLA_NET_0_74484, Y => HIEFFPLA_NET_0_74669);
    
    HIEFFPLA_INST_0_65253 : NOR3A
      port map(A => HIEFFPLA_NET_0_73430, B => 
        \Sensors_0_pressure_raw[13]\, C => 
        \Sensors_0_pressure_raw[10]\, Y => HIEFFPLA_NET_0_73434);
    
    HIEFFPLA_INST_0_66430 : NOR3B
      port map(A => HIEFFPLA_NET_0_73148, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        C => HIEFFPLA_NET_0_73043, Y => HIEFFPLA_NET_0_73123);
    
    \General_Controller_0/constant_bias_voltage_1[6]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[6]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[6]_net_1\);
    
    HIEFFPLA_INST_0_60594 : MX2
      port map(A => HIEFFPLA_NET_0_74498, B => 
        HIEFFPLA_NET_0_74428, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74390);
    
    HIEFFPLA_INST_0_65615 : NAND3
      port map(A => \Science_0/ADC_READ_0/cnt3up[3]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt3up[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt3up[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73330);
    
    HIEFFPLA_INST_0_63305 : NAND3C
      port map(A => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[4]_net_1\, C => 
        HIEFFPLA_NET_0_73810, Y => HIEFFPLA_NET_0_73782);
    
    \Science_0/ADC_READ_0/chan5_data[9]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[9]\);
    
    HIEFFPLA_INST_0_63312 : NOR3A
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        HIEFFPLA_NET_0_73786, C => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73779);
    
    HIEFFPLA_INST_0_63268 : NAND3B
      port map(A => HIEFFPLA_NET_0_73817, B => 
        HIEFFPLA_NET_0_74024, C => HIEFFPLA_NET_0_73794, Y => 
        HIEFFPLA_NET_0_73795);
    
    HIEFFPLA_INST_0_57424 : AO1
      port map(A => \Sensors_0_gyro_temp[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74874, Y => HIEFFPLA_NET_0_75050);
    
    HIEFFPLA_INST_0_64207 : MX2
      port map(A => HIEFFPLA_NET_0_73745, B => 
        HIEFFPLA_NET_0_73737, S => HIEFFPLA_NET_0_73588, Y => 
        HIEFFPLA_NET_0_73649);
    
    HIEFFPLA_INST_0_64549 : MX2A
      port map(A => HIEFFPLA_NET_0_73604, B => 
        Communications_0_uc_tx_rdy, S => HIEFFPLA_NET_0_73606, Y
         => HIEFFPLA_NET_0_73602);
    
    \General_Controller_0/status_bits_1[62]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74184, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[62]\);
    
    HIEFFPLA_INST_0_63466 : MX2
      port map(A => HIEFFPLA_NET_0_73685, B => 
        HIEFFPLA_NET_0_73677, S => HIEFFPLA_NET_0_73621, Y => 
        HIEFFPLA_NET_0_73760);
    
    \Science_0/DAC_SET_0/vector[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73193, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[3]_net_1\);
    
    HIEFFPLA_INST_0_55382 : AO1
      port map(A => HIEFFPLA_NET_0_75528, B => 
        HIEFFPLA_NET_0_75516, C => HIEFFPLA_NET_0_75513, Y => 
        HIEFFPLA_NET_0_75525);
    
    \General_Controller_0/uc_rx_byte_0[0]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[0]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte_0[0]_net_1\);
    
    HIEFFPLA_INST_0_67190 : AND3
      port map(A => HIEFFPLA_NET_0_72957, B => 
        HIEFFPLA_NET_0_72954, C => HIEFFPLA_NET_0_72952, Y => 
        HIEFFPLA_NET_0_72943);
    
    HIEFFPLA_INST_0_65135 : OA1C
      port map(A => HIEFFPLA_NET_0_73460, B => 
        HIEFFPLA_NET_0_73466, C => \Sensors_0_pressure_raw[14]\, 
        Y => HIEFFPLA_NET_0_73462);
    
    HIEFFPLA_INST_0_63758 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[5]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[5]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73716);
    
    HIEFFPLA_INST_0_60753 : MX2
      port map(A => HIEFFPLA_NET_0_74549, B => 
        HIEFFPLA_NET_0_74577, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74363);
    
    HIEFFPLA_INST_0_69708 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        C => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72324);
    
    \General_Controller_0/status_bits_1[33]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74209, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[0]\);
    
    \General_Controller_0/sweep_table_read_value[8]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74156, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[8]_net_1\);
    
    \L3WR_pad/U0/U0\ : IOPAD_TRI
      port map(D => \L3WR_pad/U0/NET1\, E => \L3WR_pad/U0/NET2\, 
        PAD => L3WR);
    
    HIEFFPLA_INST_0_62661 : AND3A
      port map(A => HIEFFPLA_NET_0_73776, B => 
        HIEFFPLA_NET_0_73860, C => HIEFFPLA_NET_0_74018, Y => 
        HIEFFPLA_NET_0_73933);
    
    HIEFFPLA_INST_0_59207 : AO1A
      port map(A => General_Controller_0_readout_en, B => 
        \GS_Readout_0/state[7]_net_1\, C => HIEFFPLA_NET_0_74582, 
        Y => HIEFFPLA_NET_0_74587);
    
    HIEFFPLA_INST_0_70252 : NOR3B
      port map(A => HIEFFPLA_NET_0_72268, B => 
        HIEFFPLA_NET_0_72284, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72186);
    
    \Timekeeper_0/microseconds[21]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72138, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[21]\);
    
    HIEFFPLA_INST_0_54931 : AX1C
      port map(A => HIEFFPLA_NET_0_75635, B => 
        HIEFFPLA_NET_0_75636, C => \ClockDivs_0/clk_800kHz_i\, Y
         => HIEFFPLA_NET_0_75637);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRY[3]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75298, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[3]\\\\\);
    
    HIEFFPLA_INST_0_67912 : AO1D
      port map(A => HIEFFPLA_NET_0_72888, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        C => HIEFFPLA_NET_0_72773, Y => HIEFFPLA_NET_0_72774);
    
    HIEFFPLA_INST_0_55128 : OA1A
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[28]_net_1\, B => 
        HIEFFPLA_NET_0_75597, C => HIEFFPLA_NET_0_75581, Y => 
        HIEFFPLA_NET_0_75582);
    
    HIEFFPLA_INST_0_70758 : AND2
      port map(A => \Timing_0/s_count[3]_net_1\, B => 
        HIEFFPLA_NET_0_72026, Y => HIEFFPLA_NET_0_72020);
    
    HIEFFPLA_INST_0_64671 : AND2
      port map(A => 
        \General_Controller_0/uc_tx_nextstate[3]_net_1\, B => 
        HIEFFPLA_NET_0_73584, Y => HIEFFPLA_NET_0_73570);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[8]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72484, Q => 
        \Sensors_0_gyro_y[8]\);
    
    HIEFFPLA_INST_0_68556 : NAND3C
      port map(A => HIEFFPLA_NET_0_72629, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, C => 
        HIEFFPLA_NET_0_72699, Y => HIEFFPLA_NET_0_72618);
    
    HIEFFPLA_INST_0_65435 : AND2B
      port map(A => \Science_0/ADC_READ_0/cnt2dn[0]_net_1\, B => 
        HIEFFPLA_NET_0_73381, Y => HIEFFPLA_NET_0_73376);
    
    HIEFFPLA_INST_0_70782 : AO1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        B => HIEFFPLA_NET_0_72013, C => HIEFFPLA_NET_0_72422, Y
         => HIEFFPLA_NET_0_72325);
    
    HIEFFPLA_INST_0_68577 : AND3A
      port map(A => HIEFFPLA_NET_0_72597, B => 
        HIEFFPLA_NET_0_72612, C => HIEFFPLA_NET_0_72623, Y => 
        HIEFFPLA_NET_0_72613);
    
    HIEFFPLA_INST_0_62780 : AND2
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73906);
    
    HIEFFPLA_INST_0_61705 : MX2
      port map(A => \SweepTable_0_RD[7]\, B => 
        \SweepTable_1_RD[7]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74157);
    
    HIEFFPLA_INST_0_60197 : MX2
      port map(A => \Science_0_chan5_data[8]\, B => 
        \Science_0_chan4_data[0]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74447);
    
    HIEFFPLA_INST_0_64705 : OR2A
      port map(A => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, B => 
        HIEFFPLA_NET_0_73552, Y => HIEFFPLA_NET_0_73558);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[10]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[10]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[10]\);
    
    HIEFFPLA_INST_0_65762 : AX1C
      port map(A => \Science_0/ADC_READ_0/cnt[3]_net_1\, B => 
        HIEFFPLA_NET_0_73297, C => 
        \Science_0/ADC_READ_0/cnt[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73286);
    
    \General_Controller_0/status_bits_1[41]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74205, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[41]\);
    
    HIEFFPLA_INST_0_63572 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[14]_net_1\, B
         => \General_Controller_0/sweep_table_points[14]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73747);
    
    HIEFFPLA_INST_0_60243 : MX2
      port map(A => HIEFFPLA_NET_0_74529, B => 
        HIEFFPLA_NET_0_74458, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74442);
    
    HIEFFPLA_INST_0_66085 : NAND2B
      port map(A => \Science_0/DAC_SET_0/state[3]_net_1\, B => 
        \Science_0/DAC_SET_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73213);
    
    HIEFFPLA_INST_0_68603 : AO1
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[5]_net_1\, B => 
        HIEFFPLA_NET_0_72705, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_72608);
    
    HIEFFPLA_INST_0_65384 : AX1C
      port map(A => \Science_0/ADC_READ_0/cnt1up[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt1up[0]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt1up[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73393);
    
    HIEFFPLA_INST_0_63734 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[1]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[1]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73720);
    
    HIEFFPLA_INST_0_56454 : XOR2
      port map(A => HIEFFPLA_NET_0_75318, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[4]\\\\\, Y => 
        HIEFFPLA_NET_0_75278);
    
    HIEFFPLA_INST_0_66568 : MX2
      port map(A => HIEFFPLA_NET_0_73089, B => 
        HIEFFPLA_NET_0_73088, S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73090);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[1]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_75252, CLK => CLKINT_0_Y_0, E
         => CLKINT_1_Y, Q => 
        \Data_Saving_0/Interrupt_Generator_0/counter[1]_net_1\);
    
    HIEFFPLA_INST_0_69617 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        B => \Sensors_0/Pressure_Sensor_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72344);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[13]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[13]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[13]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[5]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[5]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[5]\);
    
    HIEFFPLA_INST_0_69615 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72346);
    
    HIEFFPLA_INST_0_55541 : AND2
      port map(A => \Communications_0/UART_1/rx_count[2]_net_1\, 
        B => \Communications_0/UART_1/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75483);
    
    HIEFFPLA_INST_0_56042 : XA1A
      port map(A => HIEFFPLA_NET_0_75272, B => 
        HIEFFPLA_NET_0_75315, C => HIEFFPLA_NET_0_75329, Y => 
        HIEFFPLA_NET_0_75361);
    
    \Science_0/ADC_READ_0/chan7_data[10]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[10]\);
    
    HIEFFPLA_INST_0_66323 : AND2A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73146);
    
    \General_Controller_0/state_seconds[19]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74228, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[19]_net_1\);
    
    HIEFFPLA_INST_0_66900 : AO1A
      port map(A => HIEFFPLA_NET_0_73101, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        C => HIEFFPLA_NET_0_73038, Y => HIEFFPLA_NET_0_73009);
    
    HIEFFPLA_INST_0_69817 : XA1A
      port map(A => HIEFFPLA_NET_0_72303, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[4]_net_1\, 
        C => HIEFFPLA_NET_0_72236, Y => HIEFFPLA_NET_0_72296);
    
    HIEFFPLA_INST_0_55352 : NAND2
      port map(A => 
        \Communications_0/UART_0/tx_clk_count[1]_net_1\, B => 
        \Communications_0/UART_0/tx_clk_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75533);
    
    HIEFFPLA_INST_0_64520 : AO1A
      port map(A => HIEFFPLA_NET_0_73552, B => 
        HIEFFPLA_NET_0_73594, C => HIEFFPLA_NET_0_73607, Y => 
        HIEFFPLA_NET_0_73608);
    
    \Communications_0/UART_0/rx_state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75549, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/rx_state[0]_net_1\);
    
    HIEFFPLA_INST_0_56692 : MX2
      port map(A => HIEFFPLA_NET_0_75191, B => 
        HIEFFPLA_NET_0_75052, S => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75224);
    
    HIEFFPLA_INST_0_57461 : AO1
      port map(A => \Sensors_0_acc_z[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74864, Y => HIEFFPLA_NET_0_75039);
    
    HIEFFPLA_INST_0_55136 : AOI1
      port map(A => \Communications_0/UART_0/rx_clk_count_c0\, B
         => \Communications_0/UART_0/rx_clk_count[30]_net_1\, C
         => \Communications_0/UART_0/rx_clk_count[29]_net_1\, Y
         => HIEFFPLA_NET_0_75578);
    
    HIEFFPLA_INST_0_55890 : XO1A
      port map(A => HIEFFPLA_NET_0_75414, B => 
        \Communications_0/UART_1/tx_clk_count_i_0[7]\, C => 
        HIEFFPLA_NET_0_75419, Y => HIEFFPLA_NET_0_75403);
    
    HIEFFPLA_INST_0_55657 : AND2
      port map(A => \Communications_0/UART_1/rx_count[2]_net_1\, 
        B => \Communications_0/UART_1/rx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75452);
    
    \Timekeeper_0/milliseconds[21]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72103, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[21]\);
    
    HIEFFPLA_INST_0_60622 : AO1
      port map(A => HIEFFPLA_NET_0_74525, B => 
        HIEFFPLA_NET_0_74341, C => HIEFFPLA_NET_0_74505, Y => 
        HIEFFPLA_NET_0_74385);
    
    HIEFFPLA_INST_0_67777 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        B => HIEFFPLA_NET_0_72765, C => HIEFFPLA_NET_0_72903, Y
         => HIEFFPLA_NET_0_72804);
    
    HIEFFPLA_INST_0_66028 : NOR3B
      port map(A => General_Controller_0_exp_adc_reset, B => 
        HIEFFPLA_NET_0_73234, C => 
        \Science_0/ADC_RESET_0/old_enable_net_1\, Y => 
        HIEFFPLA_NET_0_73233);
    
    HIEFFPLA_INST_0_55231 : NOR2A
      port map(A => 
        \Communications_0/FFU_Command_Checker_0_rmu_oen\, B => 
        \Communications_0/UART_0/rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75556);
    
    HIEFFPLA_INST_0_70621 : XOR2
      port map(A => \Timing_0/m_time[4]_net_1\, B => 
        HIEFFPLA_NET_0_72070, Y => HIEFFPLA_NET_0_72061);
    
    HIEFFPLA_INST_0_61612 : NAND3C
      port map(A => HIEFFPLA_NET_0_74176, B => 
        HIEFFPLA_NET_0_74175, C => HIEFFPLA_NET_0_73802, Y => 
        HIEFFPLA_NET_0_74174);
    
    \General_Controller_0/constant_bias_voltage_1[7]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[7]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[7]_net_1\);
    
    \Science_0/ADC_READ_0/chan6_data[1]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[1]\);
    
    \Science_0/ADC_READ_0/chan0_data[1]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[1]\);
    
    HIEFFPLA_INST_0_63881 : AO1
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[9]_net_1\, 
        B => HIEFFPLA_NET_0_73579, C => HIEFFPLA_NET_0_73695, Y
         => HIEFFPLA_NET_0_73696);
    
    HIEFFPLA_INST_0_55512 : NOR3B
      port map(A => HIEFFPLA_NET_0_75484, B => 
        HIEFFPLA_NET_0_75488, C => 
        \Communications_0/UART_1/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75492);
    
    HIEFFPLA_INST_0_66442 : AND3C
      port map(A => HIEFFPLA_NET_0_73116, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73120);
    
    HIEFFPLA_INST_0_57283 : AND2
      port map(A => \Sensors_0_acc_y[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        Y => HIEFFPLA_NET_0_75097);
    
    HIEFFPLA_INST_0_62082 : AO1C
      port map(A => HIEFFPLA_NET_0_73875, B => 
        \General_Controller_0/uc_rx_prev_state[2]_net_1\, C => 
        HIEFFPLA_NET_0_73862, Y => HIEFFPLA_NET_0_74056);
    
    HIEFFPLA_INST_0_62123 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state_0[3]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[1]_net_1\, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74047);
    
    HIEFFPLA_INST_0_62298 : NOR3B
      port map(A => HIEFFPLA_NET_0_73970, B => 
        HIEFFPLA_NET_0_74011, C => 
        \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74012);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/num_bytes_1[1]\ : 
        DFN1
      port map(D => HIEFFPLA_NET_0_72966, CLK => CLKINT_0_Y_0, Q
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[1]\);
    
    HIEFFPLA_INST_0_70193 : AOI1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[3]_net_1\, 
        B => HIEFFPLA_NET_0_72284, C => HIEFFPLA_NET_0_72312, Y
         => HIEFFPLA_NET_0_72198);
    
    HIEFFPLA_INST_0_55344 : NAND3C
      port map(A => HIEFFPLA_NET_0_75501, B => 
        HIEFFPLA_NET_0_75533, C => 
        \Communications_0/UART_0/tx_clk_count_i_0[2]\, Y => 
        HIEFFPLA_NET_0_75536);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRYSYNC[1]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_8_Q\, CLK
         => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[1]\\\\\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[3]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72482, Q => 
        \Sensors_0_gyro_y[3]\);
    
    HIEFFPLA_INST_0_68245 : MX2A
      port map(A => HIEFFPLA_NET_0_72693, B => 
        HIEFFPLA_NET_0_72575, S => HIEFFPLA_NET_0_72622, Y => 
        HIEFFPLA_NET_0_72697);
    
    \General_Controller_0/sweep_table_read_value[2]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74162, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[2]_net_1\);
    
    \Timekeeper_0/milliseconds[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72095, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[7]\);
    
    HIEFFPLA_INST_0_56816 : MX2
      port map(A => HIEFFPLA_NET_0_75170, B => 
        HIEFFPLA_NET_0_75022, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75207);
    
    HIEFFPLA_INST_0_70390 : AND3
      port map(A => \Timekeeper_0_microseconds[9]\, B => 
        HIEFFPLA_NET_0_72157, C => 
        \Timekeeper_0_microseconds[10]\, Y => 
        HIEFFPLA_NET_0_72152);
    
    HIEFFPLA_INST_0_56865 : MX2
      port map(A => HIEFFPLA_NET_0_75005, B => 
        HIEFFPLA_NET_0_74933, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75202);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[0]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72804, Q => 
        \Sensors_0_mag_x[0]\);
    
    HIEFFPLA_INST_0_64917 : OA1C
      port map(A => HIEFFPLA_NET_0_73509, B => 
        \I2C_PassThrough_0.state[2]\, C => FRAM_SDA_in, Y => 
        HIEFFPLA_NET_0_73511);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[18]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[18]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[18]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[5]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72753, Q => 
        \Sensors_0_acc_z[5]\);
    
    HIEFFPLA_INST_0_67626 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72840);
    
    HIEFFPLA_INST_0_67223 : NAND3C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72935);
    
    HIEFFPLA_INST_0_57293 : AND2
      port map(A => \Sensors_0_gyro_x[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75087);
    
    HIEFFPLA_INST_0_56738 : AO1C
      port map(A => HIEFFPLA_NET_0_75185, B => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_75218, Y => HIEFFPLA_NET_0_75219);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[13]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72283, Q => 
        \Sensors_0_pressure_temp_raw[13]\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/state[1]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72613, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_57910 : AOI1
      port map(A => \Sensors_0_acc_time[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74907, Y => HIEFFPLA_NET_0_74908);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/data_out[3]\ : 
        DFN0E1C1
      port map(D => PRESSURE_SDA_in, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72399, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[3]\);
    
    HIEFFPLA_INST_0_65597 : XA1
      port map(A => HIEFFPLA_NET_0_73337, B => 
        \Science_0/ADC_READ_0/cnt3up[2]_net_1\, C => 
        HIEFFPLA_NET_0_73338, Y => HIEFFPLA_NET_0_73334);
    
    HIEFFPLA_INST_0_58606 : AND2B
      port map(A => \GS_Readout_0/prevState[5]_net_1\, B => 
        \GS_Readout_0/prevState[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74722);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRYSYNC[9]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_1_Q\, CLK
         => CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[9]\\\\\);
    
    HIEFFPLA_INST_0_56632 : MX2
      port map(A => HIEFFPLA_NET_0_75197, B => 
        HIEFFPLA_NET_0_75065, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75230);
    
    HIEFFPLA_INST_0_55442 : NOR3B
      port map(A => HIEFFPLA_NET_0_75510, B => 
        \Communications_0/UART_0/tx_count[0]_net_1\, C => 
        \Communications_0/UART_0/tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75512);
    
    \Science_0/ADC_READ_0/chan3_data[5]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[5]\);
    
    HIEFFPLA_INST_0_59579 : MX2
      port map(A => \Sensors_0_pressure_temp_raw[12]\, B => 
        \Sensors_0_pressure_temp_raw[16]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74535);
    
    HIEFFPLA_INST_0_67208 : XO1A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        C => HIEFFPLA_NET_0_72938, Y => HIEFFPLA_NET_0_72939);
    
    HIEFFPLA_INST_0_69069 : NOR3A
      port map(A => \Sensors_0/Gyro_0/state[8]\, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        Y => HIEFFPLA_NET_0_72478);
    
    HIEFFPLA_INST_0_68687 : OA1C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, B => 
        HIEFFPLA_NET_0_72577, C => HIEFFPLA_NET_0_72586, Y => 
        HIEFFPLA_NET_0_72587);
    
    \UC_PWR_EN_pad/U0/U0\ : IOPAD_TRI
      port map(D => \UC_PWR_EN_pad/U0/NET1\, E => 
        \UC_PWR_EN_pad/U0/NET2\, PAD => UC_PWR_EN);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[1]\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72407, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72352, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[1]_net_1\);
    
    HIEFFPLA_INST_0_60908 : AND2B
      port map(A => \General_Controller_0/un10_uc_tx_rdy_i[3]\, B
         => \General_Controller_0/un10_uc_tx_rdy_i[2]\, Y => 
        HIEFFPLA_NET_0_74322);
    
    HIEFFPLA_INST_0_63316 : NOR3A
      port map(A => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, B => 
        HIEFFPLA_NET_0_73810, C => HIEFFPLA_NET_0_73804, Y => 
        HIEFFPLA_NET_0_73778);
    
    HIEFFPLA_INST_0_58028 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_74874);
    
    HIEFFPLA_INST_0_57575 : AO1B
      port map(A => \Sensors_0_gyro_x[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75003, Y => HIEFFPLA_NET_0_75004);
    
    \GS_Readout_0/prevState[5]\ : DFN1E0C1
      port map(D => \GS_Readout_0/state[5]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \GS_Readout_0/state[6]_net_1\, Q => 
        \GS_Readout_0/prevState[5]_net_1\);
    
    \Timekeeper_0/microseconds[17]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72143, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[17]\);
    
    HIEFFPLA_INST_0_58718 : AND3
      port map(A => HIEFFPLA_NET_0_74421, B => 
        \GS_Readout_0/state[2]_net_1\, C => HIEFFPLA_NET_0_74574, 
        Y => HIEFFPLA_NET_0_74698);
    
    HIEFFPLA_INST_0_64317 : MX2
      port map(A => HIEFFPLA_NET_0_73726, B => 
        HIEFFPLA_NET_0_73718, S => HIEFFPLA_NET_0_73619, Y => 
        HIEFFPLA_NET_0_73638);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[7]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_75246, CLK => CLKINT_0_Y_0, E
         => CLKINT_1_Y, Q => 
        \Data_Saving_0/Interrupt_Generator_0/counter[7]_net_1\);
    
    HIEFFPLA_INST_0_68887 : AO1D
      port map(A => HIEFFPLA_NET_0_72514, B => 
        HIEFFPLA_NET_0_72524, C => HIEFFPLA_NET_0_72540, Y => 
        HIEFFPLA_NET_0_72532);
    
    HIEFFPLA_INST_0_62280 : AO1
      port map(A => HIEFFPLA_NET_0_74045, B => 
        HIEFFPLA_NET_0_73972, C => HIEFFPLA_NET_0_73912, Y => 
        HIEFFPLA_NET_0_74015);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72460, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\);
    
    HIEFFPLA_INST_0_57408 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_75053, Y => HIEFFPLA_NET_0_75054);
    
    HIEFFPLA_INST_0_55649 : AND2
      port map(A => HIEFFPLA_NET_0_75477, B => 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\, Y => 
        HIEFFPLA_NET_0_75455);
    
    HIEFFPLA_INST_0_58420 : NOR3A
      port map(A => \Data_Saving_0/Packet_Saver_0/mag_flag_net_1\, 
        B => \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\, C
         => \Data_Saving_0/Packet_Saver_0/acc_flag_net_1\, Y => 
        HIEFFPLA_NET_0_74772);
    
    HIEFFPLA_INST_0_62629 : NAND3C
      port map(A => HIEFFPLA_NET_0_73968, B => 
        HIEFFPLA_NET_0_73879, C => HIEFFPLA_NET_0_73957, Y => 
        HIEFFPLA_NET_0_73941);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]\ : 
        DFN0E0
      port map(D => HIEFFPLA_NET_0_73104, CLK => 
        ClockDivs_0_clk_800kHz, E => HIEFFPLA_NET_0_73056, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\);
    
    HIEFFPLA_INST_0_70615 : XOR2
      port map(A => HIEFFPLA_NET_0_72068, B => 
        \Timing_0/m_time[6]_net_1\, Y => HIEFFPLA_NET_0_72063);
    
    HIEFFPLA_INST_0_56534 : AX1C
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[3]_net_1\, B
         => HIEFFPLA_NET_0_75256, C => 
        \Data_Saving_0/Interrupt_Generator_0/counter[4]_net_1\, Y
         => HIEFFPLA_NET_0_75249);
    
    \FRAM_SCL_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => FRAM_SCL_c_c, E => \VCC\, DOUT => 
        \FRAM_SCL_pad/U0/NET1\, EOUT => \FRAM_SCL_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_58927 : NOR3B
      port map(A => HIEFFPLA_NET_0_74359, B => 
        HIEFFPLA_NET_0_74649, C => HIEFFPLA_NET_0_74421, Y => 
        HIEFFPLA_NET_0_74657);
    
    \General_Controller_0/constant_bias_voltage_1[8]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[8]_net_1\);
    
    HIEFFPLA_INST_0_57355 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_74855, Y => HIEFFPLA_NET_0_75068);
    
    HIEFFPLA_INST_0_70104 : AOI1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[2]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        C => HIEFFPLA_NET_0_72271, Y => HIEFFPLA_NET_0_72218);
    
    HIEFFPLA_INST_0_59321 : NOR3B
      port map(A => HIEFFPLA_NET_0_74433, B => 
        HIEFFPLA_NET_0_74405, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74569);
    
    \General_Controller_0/uc_rx_byte[5]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[5]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte[5]_net_1\);
    
    HIEFFPLA_INST_0_60344 : MX2
      port map(A => HIEFFPLA_NET_0_74460, B => 
        HIEFFPLA_NET_0_74512, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74429);
    
    HIEFFPLA_INST_0_64151 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_1[4]_net_1\, 
        B => 
        \General_Controller_0/constant_bias_voltage_1[12]_net_1\, 
        S => \General_Controller_0/uc_tx_substate[1]_net_1\, Y
         => HIEFFPLA_NET_0_73661);
    
    HIEFFPLA_INST_0_67016 : NOR3A
      port map(A => HIEFFPLA_NET_0_72976, B => 
        HIEFFPLA_NET_0_72890, C => HIEFFPLA_NET_0_72913, Y => 
        HIEFFPLA_NET_0_72984);
    
    HIEFFPLA_INST_0_66253 : XO1
      port map(A => \Science_0/SET_LP_GAIN_0/old_G4[1]_net_1\, B
         => \Science_0/ADC_READ_0_G4[1]\, C => 
        HIEFFPLA_NET_0_73165, Y => HIEFFPLA_NET_0_73166);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[11]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[11]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[11]\);
    
    HIEFFPLA_INST_0_64010 : MX2
      port map(A => HIEFFPLA_NET_0_73651, B => 
        HIEFFPLA_NET_0_73643, S => HIEFFPLA_NET_0_73599, Y => 
        HIEFFPLA_NET_0_73680);
    
    HIEFFPLA_INST_0_61171 : NAND3C
      port map(A => HIEFFPLA_NET_0_74258, B => 
        \General_Controller_0/state_seconds[15]_net_1\, C => 
        HIEFFPLA_NET_0_74242, Y => HIEFFPLA_NET_0_74259);
    
    \Communications_0/UART_0/recv[3]\ : DFN1E1C1
      port map(D => \Communications_0/UART_0/rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75551, Q => 
        \Communications_0/UART_0_recv[3]\);
    
    HIEFFPLA_INST_0_70063 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]_net_1\, 
        B => HIEFFPLA_NET_0_72237, C => HIEFFPLA_NET_0_72226, Y
         => HIEFFPLA_NET_0_72231);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[3]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73136, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[3]_net_1\);
    
    HIEFFPLA_INST_0_68984 : AND3C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[5]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[6]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72507);
    
    HIEFFPLA_INST_0_69899 : NAND2B
      port map(A => HIEFFPLA_NET_0_72278, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72273);
    
    \Science_0/ADC_READ_0/cnt_chan[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73279, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/ADC_READ_0/cnt_chan[0]_net_1\);
    
    HIEFFPLA_INST_0_60268 : MX2
      port map(A => HIEFFPLA_NET_0_74362, B => 
        HIEFFPLA_NET_0_74388, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74439);
    
    HIEFFPLA_INST_0_70472 : AND3
      port map(A => \Timekeeper_0_milliseconds[9]\, B => 
        HIEFFPLA_NET_0_72124, C => 
        \Timekeeper_0_milliseconds[10]\, Y => 
        HIEFFPLA_NET_0_72119);
    
    HIEFFPLA_INST_0_66720 : AO1A
      port map(A => HIEFFPLA_NET_0_73113, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_73055);
    
    HIEFFPLA_INST_0_58207 : AO1
      port map(A => \ch3_data_net_0[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74828, Y => HIEFFPLA_NET_0_74829);
    
    HIEFFPLA_INST_0_69289 : OR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72429);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72472, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]_net_1\);
    
    HIEFFPLA_INST_0_58435 : NOR3B
      port map(A => HIEFFPLA_NET_0_74771, B => 
        \Data_Saving_0/Packet_Saver_0/pressure_flag_net_1\, C => 
        \Data_Saving_0/Packet_Saver_0/gyro_flag_net_1\, Y => 
        HIEFFPLA_NET_0_74767);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[15]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[15]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[15]\);
    
    HIEFFPLA_INST_0_59627 : MX2
      port map(A => \Science_0_chan1_data[0]\, B => 
        \Science_0_chan1_data[4]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74529);
    
    HIEFFPLA_INST_0_68215 : AO1A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\, B => 
        HIEFFPLA_NET_0_72702, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, Y => 
        HIEFFPLA_NET_0_72704);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_RNIRAS8[9]\ : 
        CLKINT
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[9]\, Y => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\);
    
    \Communications_0/UART_1/rx_clk_count[29]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75458, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75443, Q => 
        \Communications_0/UART_1/rx_clk_count[29]_net_1\);
    
    HIEFFPLA_INST_0_62830 : OA1C
      port map(A => HIEFFPLA_NET_0_73940, B => 
        HIEFFPLA_NET_0_73810, C => HIEFFPLA_NET_0_73910, Y => 
        HIEFFPLA_NET_0_73891);
    
    \Science_0/ADC_READ_0/chan7_data[1]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[1]\);
    
    HIEFFPLA_INST_0_68707 : NOR2A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\, B
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0_we\, Y => 
        HIEFFPLA_NET_0_72582);
    
    HIEFFPLA_INST_0_58454 : AXO2
      port map(A => \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, 
        B => General_Controller_0_en_data_saving, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74762);
    
    HIEFFPLA_INST_0_57322 : AO1
      port map(A => \Sensors_0_gyro_z[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75076, Y => HIEFFPLA_NET_0_75077);
    
    HIEFFPLA_INST_0_70271 : AO1
      port map(A => HIEFFPLA_NET_0_72176, B => 
        HIEFFPLA_NET_0_72175, C => HIEFFPLA_NET_0_72202, Y => 
        HIEFFPLA_NET_0_72182);
    
    HIEFFPLA_INST_0_69443 : AND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72388);
    
    HIEFFPLA_INST_0_64662 : NOR3B
      port map(A => HIEFFPLA_NET_0_73920, B => 
        HIEFFPLA_NET_0_73565, C => HIEFFPLA_NET_0_73584, Y => 
        HIEFFPLA_NET_0_73573);
    
    \General_Controller_0/sweep_table_write_value[11]\ : DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[11]_net_1\);
    
    \Timing_0/f_time[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72086, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \s_clks_net_0[4]\);
    
    HIEFFPLA_INST_0_70967 : MX2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[1]\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[3]\, 
        S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72000);
    
    HIEFFPLA_INST_0_64515 : NOR2A
      port map(A => HIEFFPLA_NET_0_73617, B => 
        HIEFFPLA_NET_0_73933, Y => HIEFFPLA_NET_0_73609);
    
    HIEFFPLA_INST_0_55373 : AOI1C
      port map(A => \Communications_0/UART_0/tx_state[0]_net_1\, 
        B => \Communications_0/UART_0/tx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_75528, Y => HIEFFPLA_NET_0_75527);
    
    HIEFFPLA_INST_0_62653 : AND3C
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[1]_net_1\, C => 
        HIEFFPLA_NET_0_73935, Y => HIEFFPLA_NET_0_73936);
    
    HIEFFPLA_INST_0_55174 : XA1B
      port map(A => \Communications_0/UART_0/rx_clk_count_c0\, B
         => \Communications_0/UART_0/rx_clk_count[30]_net_1\, C
         => HIEFFPLA_NET_0_75567, Y => HIEFFPLA_NET_0_75569);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_WRITE_RESET_P_0\ : DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_12_Q\, 
        CLK => CLKINT_0_Y_0, CLR => \AFLSDF_INV_12\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\);
    
    HIEFFPLA_INST_0_68073 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, Y
         => HIEFFPLA_NET_0_72740);
    
    HIEFFPLA_INST_0_65377 : NOR3B
      port map(A => HIEFFPLA_NET_0_73276, B => 
        HIEFFPLA_NET_0_73395, C => 
        \Science_0/ADC_READ_0/cnt1up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73396);
    
    HIEFFPLA_INST_0_57416 : AO1
      port map(A => \Sensors_0_gyro_temp[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75051, Y => HIEFFPLA_NET_0_75052);
    
    HIEFFPLA_INST_0_63275 : AND2
      port map(A => \General_Controller_0/uc_rx_state_0[1]_net_1\, 
        B => \General_Controller_0/uc_rx_substate[0]_net_1\, Y
         => HIEFFPLA_NET_0_73793);
    
    HIEFFPLA_INST_0_57257 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[51]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75107);
    
    HIEFFPLA_INST_0_69905 : OR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        C => HIEFFPLA_NET_0_72267, Y => HIEFFPLA_NET_0_72270);
    
    HIEFFPLA_INST_0_65348 : XA1B
      port map(A => HIEFFPLA_NET_0_73413, B => 
        \Science_0/ADC_READ_0/cnt1dn[5]_net_1\, C => 
        HIEFFPLA_NET_0_73244, Y => HIEFFPLA_NET_0_73403);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[19]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72280, Q => \Sensors_0_pressure_raw[19]\);
    
    HIEFFPLA_INST_0_61772 : AX1C
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[13]_net_1\, B
         => HIEFFPLA_NET_0_74147, C => 
        \General_Controller_0/sweep_table_sweep_cnt[14]_net_1\, Y
         => HIEFFPLA_NET_0_74139);
    
    HIEFFPLA_INST_0_58270 : AO1
      port map(A => \Sensors_0_mag_x[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_75123, Y => HIEFFPLA_NET_0_74815);
    
    HIEFFPLA_INST_0_59441 : MX2
      port map(A => HIEFFPLA_NET_0_74396, B => 
        HIEFFPLA_NET_0_74464, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74554);
    
    HIEFFPLA_INST_0_65624 : AND2
      port map(A => HIEFFPLA_NET_0_73329, B => 
        \Science_0/ADC_READ_0/cnt4dn[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73326);
    
    \General_Controller_0/uc_rx_substate[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73772, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_substate[2]_net_1\);
    
    \Eject_Signal_Debounce_0/ms_cnt[5]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74741, CLK => CLKINT_0_Y_0, Q
         => \Eject_Signal_Debounce_0/ms_cnt[5]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_1[5]\ : DFN0E0C1
      port map(D => 
        \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\);
    
    HIEFFPLA_INST_0_55949 : AXOI7
      port map(A => \Communications_0/UART_1/tx_state[0]_net_1\, 
        B => \Communications_0/UART_1/tx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_75420, Y => HIEFFPLA_NET_0_75387);
    
    HIEFFPLA_INST_0_70565 : AX1C
      port map(A => \Timing_0/m_count[0]_net_1\, B => 
        \Timing_0/m_count[1]_net_1\, C => 
        \Timing_0/m_count[2]_net_1\, Y => HIEFFPLA_NET_0_72078);
    
    HIEFFPLA_INST_0_57215 : AND2
      port map(A => \Sensors_0_acc_time[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, Y
         => HIEFFPLA_NET_0_75126);
    
    HIEFFPLA_INST_0_67496 : AO1D
      port map(A => HIEFFPLA_NET_0_72852, B => 
        HIEFFPLA_NET_0_72833, C => HIEFFPLA_NET_0_72937, Y => 
        HIEFFPLA_NET_0_72865);
    
    HIEFFPLA_INST_0_65430 : NAND2B
      port map(A => \Science_0/ADC_READ_0/cnt2dn[4]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2dn[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73378);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_10\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[0]\\\\\, CLK => 
        CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_10_Q\);
    
    HIEFFPLA_INST_0_68659 : AND3
      port map(A => HIEFFPLA_NET_0_72689, B => 
        HIEFFPLA_NET_0_72583, C => HIEFFPLA_NET_0_72662, Y => 
        HIEFFPLA_NET_0_72595);
    
    HIEFFPLA_INST_0_57330 : AO1B
      port map(A => \Sensors_0_gyro_z[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75074, Y => HIEFFPLA_NET_0_75075);
    
    HIEFFPLA_INST_0_70447 : AND3
      port map(A => \Timekeeper_0_milliseconds[19]\, B => 
        HIEFFPLA_NET_0_72123, C => 
        \Timekeeper_0_milliseconds[20]\, Y => 
        HIEFFPLA_NET_0_72126);
    
    HIEFFPLA_INST_0_62439 : NAND3C
      port map(A => \General_Controller_0/uc_rx_state_0[4]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[0]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73982);
    
    HIEFFPLA_INST_0_71053 : AO1
      port map(A => \General_Controller_0/uc_rx_byte[0]_net_1\, B
         => HIEFFPLA_NET_0_74080, C => HIEFFPLA_NET_0_71985, Y
         => HIEFFPLA_NET_0_73819);
    
    HIEFFPLA_INST_0_69546 : MX2
      port map(A => HIEFFPLA_NET_0_72344, B => 
        \Sensors_0.Pressure_Sensor_0.I2C_Master_0.sda_1\, S => 
        HIEFFPLA_NET_0_72376, Y => HIEFFPLA_NET_0_72367);
    
    HIEFFPLA_INST_0_60735 : MX2
      port map(A => \Science_0_chan2_data[7]\, B => 
        \Science_0_chan2_data[11]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74366);
    
    \General_Controller_0/constant_bias_voltage_1[3]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[3]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[3]_net_1\);
    
    HIEFFPLA_INST_0_58603 : NOR3A
      port map(A => \GS_Readout_0/state[6]_net_1\, B => 
        \GS_Readout_0/prevState[1]_net_1\, C => 
        Communications_0_ext_tx_rdy, Y => HIEFFPLA_NET_0_74724);
    
    HIEFFPLA_INST_0_61258 : XA1C
      port map(A => 
        \General_Controller_0/state_seconds[14]_net_1\, B => 
        HIEFFPLA_NET_0_74244, C => HIEFFPLA_NET_0_74217, Y => 
        HIEFFPLA_NET_0_74235);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[20]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[20]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[20]\);
    
    HIEFFPLA_INST_0_58358 : AO1
      port map(A => \Sensors_0_mag_y[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75104, Y => HIEFFPLA_NET_0_74793);
    
    AFLSDF_INV_23 : INV
      port map(A => Science_0_exp_new_data, Y => \AFLSDF_INV_23\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[21]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[21]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[21]\);
    
    HIEFFPLA_INST_0_55122 : AO1C
      port map(A => HIEFFPLA_NET_0_75587, B => 
        HIEFFPLA_NET_0_75585, C => 
        \Communications_0/UART_0/rx_clk_count[23]_net_1\, Y => 
        HIEFFPLA_NET_0_75583);
    
    HIEFFPLA_INST_0_67324 : NOR3A
      port map(A => HIEFFPLA_NET_0_72908, B => 
        HIEFFPLA_NET_0_72739, C => HIEFFPLA_NET_0_72799, Y => 
        HIEFFPLA_NET_0_72907);
    
    HIEFFPLA_INST_0_66533 : AO1
      port map(A => HIEFFPLA_NET_0_73059, B => ACCE_SCL_c, C => 
        HIEFFPLA_NET_0_73047, Y => HIEFFPLA_NET_0_73100);
    
    HIEFFPLA_INST_0_58561 : MX2
      port map(A => \Eject_Signal_Debounce_0/state[1]_net_1\, B
         => FFU_EJECTED_c, S => HIEFFPLA_NET_0_74749, Y => 
        HIEFFPLA_NET_0_74734);
    
    HIEFFPLA_INST_0_56351 : XNOR3
      port map(A => HIEFFPLA_NET_0_75265, B => 
        HIEFFPLA_NET_0_75350, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, Y
         => HIEFFPLA_NET_0_75303);
    
    \General_Controller_0/st_waddr[1]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[1]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_waddr[1]\);
    
    HIEFFPLA_INST_0_70529 : AX1C
      port map(A => \Timekeeper_0_milliseconds[7]\, B => 
        HIEFFPLA_NET_0_72120, C => \Timekeeper_0_milliseconds[8]\, 
        Y => HIEFFPLA_NET_0_72094);
    
    HIEFFPLA_INST_0_69101 : NAND3C
      port map(A => HIEFFPLA_NET_0_72458, B => 
        HIEFFPLA_NET_0_72499, C => HIEFFPLA_NET_0_72452, Y => 
        HIEFFPLA_NET_0_72470);
    
    HIEFFPLA_INST_0_55861 : AO1
      port map(A => HIEFFPLA_NET_0_75420, B => 
        HIEFFPLA_NET_0_75401, C => HIEFFPLA_NET_0_75397, Y => 
        HIEFFPLA_NET_0_75410);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRYSYNC[6]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_15_Q\, 
        CLK => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[6]\\\\\);
    
    HIEFFPLA_INST_0_65852 : MX2
      port map(A => \Science_0/ADC_READ_0_G1[0]\, B => 
        \Science_0/ADC_READ_0_G3[0]\, S => 
        \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73270);
    
    HIEFFPLA_INST_0_56057 : XA1A
      port map(A => HIEFFPLA_NET_0_75265, B => 
        HIEFFPLA_NET_0_75271, C => HIEFFPLA_NET_0_75357, Y => 
        HIEFFPLA_NET_0_75358);
    
    HIEFFPLA_INST_0_58530 : AO1
      port map(A => HIEFFPLA_NET_0_74731, B => 
        HIEFFPLA_NET_0_74738, C => HIEFFPLA_NET_0_74740, Y => 
        HIEFFPLA_NET_0_74742);
    
    HIEFFPLA_INST_0_57943 : AO1
      port map(A => \Science_0_exp_packet_0[69]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75164, Y => HIEFFPLA_NET_0_74898);
    
    HIEFFPLA_INST_0_69193 : AND3B
      port map(A => HIEFFPLA_NET_0_72439, B => 
        HIEFFPLA_NET_0_72487, C => HIEFFPLA_NET_0_72505, Y => 
        HIEFFPLA_NET_0_72450);
    
    HIEFFPLA_INST_0_65575 : XA1
      port map(A => HIEFFPLA_NET_0_73339, B => 
        \Science_0/ADC_READ_0/cnt3dn[7]_net_1\, C => 
        HIEFFPLA_NET_0_73349, Y => HIEFFPLA_NET_0_73340);
    
    \Science_0/ADC_READ_0/chan4_data[7]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[7]\);
    
    HIEFFPLA_INST_0_68513 : AO1
      port map(A => HIEFFPLA_NET_0_72620, B => GYRO_SCL_c, C => 
        \Sensors_0/Gyro_0/state[8]\, Y => HIEFFPLA_NET_0_72632);
    
    HIEFFPLA_INST_0_54949 : AX1C
      port map(A => \ClockDivs_0/cnt_800kHz[3]_net_1\, B => 
        HIEFFPLA_NET_0_75632, C => 
        \ClockDivs_0/cnt_800kHz[4]_net_1\, Y => 
        HIEFFPLA_NET_0_75631);
    
    AFLSDF_INV_14 : INV
      port map(A => \s_clks_net_0[18]\, Y => \AFLSDF_INV_14\);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_DVLDI\ : DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/MEMRENEG\, CLK
         => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\);
    
    HIEFFPLA_INST_0_59653 : MX2
      port map(A => HIEFFPLA_NET_0_74502, B => 
        HIEFFPLA_NET_0_74557, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74526);
    
    \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[1]\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72687, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72618, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[1]_net_1\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/data_out[2]\ : 
        DFN0E1C1
      port map(D => ACCE_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73123, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\);
    
    HIEFFPLA_INST_0_68835 : NOR3B
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, C
         => CLKINT_1_Y, Y => HIEFFPLA_NET_0_72545);
    
    \General_Controller_0/sweep_table_sample_skip[4]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[4]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[4]_net_1\);
    
    HIEFFPLA_INST_0_62688 : AND3B
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => HIEFFPLA_NET_0_73875, C => HIEFFPLA_NET_0_73937, Y
         => HIEFFPLA_NET_0_73928);
    
    HIEFFPLA_INST_0_61283 : XA1C
      port map(A => 
        \General_Controller_0/state_seconds[19]_net_1\, B => 
        HIEFFPLA_NET_0_74215, C => HIEFFPLA_NET_0_74217, Y => 
        HIEFFPLA_NET_0_74228);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/temp[2]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72907, Q => 
        \Sensors_0_acc_temp[2]\);
    
    HIEFFPLA_INST_0_66294 : AO1C
      port map(A => HIEFFPLA_NET_0_73179, B => 
        \Science_0/SET_LP_GAIN_0/state[7]_net_1\, C => 
        \Science_0/SET_LP_GAIN_0/state_i_0[3]\, Y => 
        HIEFFPLA_NET_0_73153);
    
    HIEFFPLA_INST_0_64397 : MX2
      port map(A => HIEFFPLA_NET_0_73710, B => 
        HIEFFPLA_NET_0_73702, S => HIEFFPLA_NET_0_73593, Y => 
        HIEFFPLA_NET_0_73630);
    
    \FMC_DA_pad[4]/U0/U0\ : IOPAD_TRI
      port map(D => \FMC_DA_pad[4]/U0/NET1\, E => 
        \FMC_DA_pad[4]/U0/NET2\, PAD => FMC_DA(4));
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[7]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72276, Q => \Sensors_0_pressure_raw[7]\);
    
    HIEFFPLA_INST_0_63752 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[4]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[4]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73717);
    
    \Science_0/ADC_READ_0/chan1_data[4]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[4]\);
    
    HIEFFPLA_INST_0_55984 : MX2
      port map(A => \Communications_0/UART_1_tx\, B => 
        HIEFFPLA_NET_0_75638, S => UC_CONSOLE_EN_c, Y => 
        UC_UART_RX_c);
    
    HIEFFPLA_INST_0_55895 : AO1
      port map(A => HIEFFPLA_NET_0_75398, B => 
        \Communications_0/UART_1/tx_clk_count_i_0[8]\, C => 
        HIEFFPLA_NET_0_75419, Y => HIEFFPLA_NET_0_75402);
    
    HIEFFPLA_INST_0_55805 : MX2C
      port map(A => \Communications_0/UART_1/tx_byte[2]_net_1\, B
         => \Communications_0/UART_1/tx_byte[6]_net_1\, S => 
        \Communications_0/UART_1/tx_count[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75423);
    
    HIEFFPLA_INST_0_88378 : AO1B
      port map(A => HIEFFPLA_NET_0_75341, B => 
        HIEFFPLA_NET_0_75336, C => HIEFFPLA_NET_0_88380, Y => 
        HIEFFPLA_NET_0_88381);
    
    AFLSDF_INV_26 : INV
      port map(A => \s_clks_net_0[9]\, Y => \AFLSDF_INV_26\);
    
    HIEFFPLA_INST_0_64879 : NOR3B
      port map(A => \I2C_PassThrough_0/cnt[4]_net_1\, B => 
        \I2C_PassThrough_0/cnt[2]_net_1\, C => 
        \I2C_PassThrough_0/cnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73519);
    
    HIEFFPLA_INST_0_57539 : AO1B
      port map(A => \Sensors_0_gyro_z[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75015, Y => HIEFFPLA_NET_0_75016);
    
    HIEFFPLA_INST_0_67669 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, B
         => \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72828);
    
    HIEFFPLA_INST_0_68162 : AO1D
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => \Sensors_0/Accelerometer_0/state[8]\, C => 
        HIEFFPLA_NET_0_72718, Y => HIEFFPLA_NET_0_72719);
    
    HIEFFPLA_INST_0_59204 : NAND3B
      port map(A => HIEFFPLA_NET_0_74360, B => 
        HIEFFPLA_NET_0_74387, C => \GS_Readout_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_74588);
    
    HIEFFPLA_INST_0_58032 : AO1
      port map(A => \Sensors_0_mag_y[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75162, Y => HIEFFPLA_NET_0_74872);
    
    HIEFFPLA_INST_0_66681 : NOR3B
      port map(A => HIEFFPLA_NET_0_73046, B => 
        HIEFFPLA_NET_0_73065, C => HIEFFPLA_NET_0_73132, Y => 
        HIEFFPLA_NET_0_73066);
    
    HIEFFPLA_INST_0_60959 : NAND2B
      port map(A => \Timekeeper_0_milliseconds[8]\, B => 
        HIEFFPLA_NET_0_74281, Y => HIEFFPLA_NET_0_74310);
    
    \General_Controller_0/sweep_table_samples_per_point[3]\ : 
        DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[3]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[3]_net_1\);
    
    HIEFFPLA_INST_0_65912 : OA1A
      port map(A => HIEFFPLA_NET_0_73365, B => 
        \Science_0/ADC_READ_0_G2[1]\, C => HIEFFPLA_NET_0_73382, 
        Y => HIEFFPLA_NET_0_73259);
    
    HIEFFPLA_INST_0_56501 : AX1C
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, B
         => HIEFFPLA_NET_0_75351, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\, Y
         => HIEFFPLA_NET_0_75262);
    
    \General_Controller_0/sweep_table_sweep_cnt[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74131, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[7]_net_1\);
    
    \Communications_0/UART_1/rx_count[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75449, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75442, Q => 
        \Communications_0/UART_1/rx_count[1]_net_1\);
    
    HIEFFPLA_INST_0_60982 : MX2A
      port map(A => General_Controller_0_exp_adc_reset, B => 
        HIEFFPLA_NET_0_74249, S => HIEFFPLA_NET_0_74339, Y => 
        HIEFFPLA_NET_0_74304);
    
    \Science_0/ADC_READ_0/exp_packet_1[36]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[2]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[36]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[17]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[1]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[17]\);
    
    HIEFFPLA_INST_0_57400 : AO1
      port map(A => \Sensors_0_gyro_temp[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75055, Y => HIEFFPLA_NET_0_75056);
    
    HIEFFPLA_INST_0_57368 : AO1
      port map(A => \ch3_data_net_0[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75064, Y => HIEFFPLA_NET_0_75065);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[1]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72279, Q => 
        \Sensors_0_pressure_temp_raw[1]\);
    
    HIEFFPLA_INST_0_55966 : AO1
      port map(A => \Communications_0/UART_1/tx_state[0]_net_1\, 
        B => HIEFFPLA_NET_0_75420, C => HIEFFPLA_NET_0_75381, Y
         => HIEFFPLA_NET_0_75382);
    
    \General_Controller_0/temp_first_byte[0]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73872, Q => 
        \General_Controller_0/temp_first_byte[0]_net_1\);
    
    HIEFFPLA_INST_0_60842 : AND3
      port map(A => HIEFFPLA_NET_0_74345, B => 
        \GS_Readout_0/subState[2]_net_1\, C => 
        \GS_Readout_0/subState[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74347);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[10]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72553, Q => 
        \Sensors_0_gyro_x[10]\);
    
    HIEFFPLA_INST_0_68425 : NAND2B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[1]\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72653);
    
    HIEFFPLA_INST_0_62893 : OR3A
      port map(A => \General_Controller_0/uc_rx_state[3]_net_1\, 
        B => HIEFFPLA_NET_0_73785, C => 
        \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73873);
    
    HIEFFPLA_INST_0_58843 : NOR3B
      port map(A => HIEFFPLA_NET_0_74490, B => 
        HIEFFPLA_NET_0_74646, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74675);
    
    HIEFFPLA_INST_0_58020 : AOI1
      port map(A => \Sensors_0_acc_time[17]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74876, Y => HIEFFPLA_NET_0_74877);
    
    HIEFFPLA_INST_0_57907 : AO1B
      port map(A => \Sensors_0_mag_time[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74908, Y => HIEFFPLA_NET_0_74909);
    
    HIEFFPLA_INST_0_56722 : MX2
      port map(A => HIEFFPLA_NET_0_75188, B => 
        HIEFFPLA_NET_0_75048, S => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75221);
    
    HIEFFPLA_INST_0_69869 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72284);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[1]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72754, Q => 
        \Sensors_0_acc_z[1]\);
    
    HIEFFPLA_INST_0_61934 : NOR3A
      port map(A => HIEFFPLA_NET_0_74022, B => 
        HIEFFPLA_NET_0_73799, C => HIEFFPLA_NET_0_74114, Y => 
        HIEFFPLA_NET_0_74095);
    
    HIEFFPLA_INST_0_70107 : NOR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        B => HIEFFPLA_NET_0_72240, C => HIEFFPLA_NET_0_72269, Y
         => HIEFFPLA_NET_0_72217);
    
    HIEFFPLA_INST_0_62758 : AO1A
      port map(A => HIEFFPLA_NET_0_73944, B => 
        HIEFFPLA_NET_0_73943, C => HIEFFPLA_NET_0_73911, Y => 
        HIEFFPLA_NET_0_73912);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[19]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[19]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[19]\);
    
    HIEFFPLA_INST_0_65241 : NOR3B
      port map(A => HIEFFPLA_NET_0_73435, B => 
        HIEFFPLA_NET_0_73429, C => HIEFFPLA_NET_0_73427, Y => 
        HIEFFPLA_NET_0_73436);
    
    HIEFFPLA_INST_0_55062 : NOR2A
      port map(A => \Communications_0/UART_0/rx_count[2]_net_1\, 
        B => \Communications_0/UART_0/rx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75600);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[23]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[23]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[23]\);
    
    HIEFFPLA_INST_0_69672 : OA1C
      port map(A => HIEFFPLA_NET_0_72382, B => 
        HIEFFPLA_NET_0_72344, C => HIEFFPLA_NET_0_72328, Y => 
        HIEFFPLA_NET_0_72332);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[5]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72276, Q => \Sensors_0_pressure_raw[5]\);
    
    HIEFFPLA_INST_0_62325 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state_0[3]_net_1\, 
        B => HIEFFPLA_NET_0_73908, C => 
        \General_Controller_0/uc_rx_state_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74005);
    
    \General_Controller_0/sweep_table_sample_skip[7]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[7]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[7]_net_1\);
    
    \Timing_0/f_time[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72089, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/f_time[1]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[3]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72754, Q => 
        \Sensors_0_acc_z[3]\);
    
    \Data_Saving_0/Packet_Saver_0/data_out[6]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75207, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[6]\);
    
    HIEFFPLA_INST_0_70095 : AND2
      port map(A => \Eject_Signal_Debounce_0/old_1kHz_i_0\, B => 
        \m_time[7]\, Y => HIEFFPLA_NET_0_72220);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72769, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\);
    
    \Communications_0/UART_0/tx_clk_count[4]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75522, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_clk_count_i_0[4]\);
    
    HIEFFPLA_INST_0_55954 : AND2B
      port map(A => \Communications_0/UART_1/tx_state[0]_net_1\, 
        B => \Communications_0/UART_1/tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75386);
    
    HIEFFPLA_INST_0_68474 : AOI1A
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, C
         => HIEFFPLA_NET_0_72641, Y => HIEFFPLA_NET_0_72642);
    
    HIEFFPLA_INST_0_66733 : NOR3B
      port map(A => HIEFFPLA_NET_0_73144, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        C => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73051);
    
    HIEFFPLA_INST_0_70312 : NOR3B
      port map(A => HIEFFPLA_NET_0_72196, B => 
        HIEFFPLA_NET_0_72195, C => HIEFFPLA_NET_0_72285, Y => 
        HIEFFPLA_NET_0_72176);
    
    HIEFFPLA_INST_0_69614 : AND3
      port map(A => PRESSURE_SCL_c, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        C => PRESSURE_SDA_in, Y => HIEFFPLA_NET_0_72347);
    
    HIEFFPLA_INST_0_66867 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_repeat_start\, 
        Y => HIEFFPLA_NET_0_73017);
    
    \General_Controller_0/sweep_table_samples_per_step[2]\ : 
        DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[2]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[2]_net_1\);
    
    HIEFFPLA_INST_0_71008 : AND3A
      port map(A => HIEFFPLA_NET_0_71991, B => 
        \Pressure_Signal_Debounce_0/ms_cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_73478, Y => HIEFFPLA_NET_0_73444);
    
    HIEFFPLA_INST_0_67439 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, Y
         => HIEFFPLA_NET_0_72880);
    
    HIEFFPLA_INST_0_61516 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[57]\, B => 
        \Timekeeper_0_milliseconds[17]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74189);
    
    HIEFFPLA_INST_0_57088 : NAND3B
      port map(A => HIEFFPLA_NET_0_74870, B => 
        HIEFFPLA_NET_0_74871, C => HIEFFPLA_NET_0_75169, Y => 
        HIEFFPLA_NET_0_75170);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[14]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[14]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[14]\);
    
    HIEFFPLA_INST_0_60897 : AND3C
      port map(A => \General_Controller_0/command[2]_net_1\, B
         => \General_Controller_0/command[1]_net_1\, C => 
        \General_Controller_0/command[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74326);
    
    HIEFFPLA_INST_0_58477 : NOR2A
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/status_flag_net_1\, B => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74757);
    
    \GS_Readout_0/subState[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74353, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/subState[2]_net_1\);
    
    HIEFFPLA_INST_0_63584 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[8]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_sample_skip[8]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73745);
    
    \Communications_0/UART_1/tx\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75428, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => \Communications_0/UART_1_tx\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[12]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[12]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[12]\);
    
    HIEFFPLA_INST_0_55632 : XA1
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[27]_net_1\, B => 
        HIEFFPLA_NET_0_75454, C => HIEFFPLA_NET_0_75437, Y => 
        HIEFFPLA_NET_0_75460);
    
    HIEFFPLA_INST_0_69822 : XA1
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[5]_net_1\, 
        B => HIEFFPLA_NET_0_72294, C => HIEFFPLA_NET_0_72236, Y
         => HIEFFPLA_NET_0_72295);
    
    HIEFFPLA_INST_0_55870 : XO1A
      port map(A => HIEFFPLA_NET_0_75418, B => 
        \Communications_0/UART_1/tx_clk_count_i_0[3]\, C => 
        HIEFFPLA_NET_0_75419, Y => HIEFFPLA_NET_0_75408);
    
    HIEFFPLA_INST_0_65550 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt3dn[2]_net_1\, B => 
        HIEFFPLA_NET_0_73354, C => HIEFFPLA_NET_0_73349, Y => 
        HIEFFPLA_NET_0_73345);
    
    \General_Controller_0/uc_rx_substate[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73773, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_substate[1]_net_1\);
    
    HIEFFPLA_INST_0_65458 : XA1C
      port map(A => \Science_0/ADC_READ_0/cnt2dn[5]_net_1\, B => 
        HIEFFPLA_NET_0_73379, C => HIEFFPLA_NET_0_73381, Y => 
        HIEFFPLA_NET_0_73371);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[11]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[11]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[11]\);
    
    HIEFFPLA_INST_0_70736 : XOR2
      port map(A => \Timing_0/m_count[0]_net_1\, B => 
        \Timing_0/m_count[1]_net_1\, Y => HIEFFPLA_NET_0_72027);
    
    HIEFFPLA_INST_0_64173 : AOI1C
      port map(A => \General_Controller_0/uc_tx_state[14]_net_1\, 
        B => HIEFFPLA_NET_0_73753, C => 
        \General_Controller_0/uc_tx_state[12]_net_1\, Y => 
        HIEFFPLA_NET_0_73657);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]\ : 
        DFN0E0
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        CLK => ClockDivs_0_clk_800kHz, E => HIEFFPLA_NET_0_73056, 
        Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\);
    
    \Science_0/ADC_READ_0/cnt1dn[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73407, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1dn[1]_net_1\);
    
    HIEFFPLA_INST_0_57389 : AND2
      port map(A => \Science_0_exp_packet_0[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        Y => HIEFFPLA_NET_0_75059);
    
    \Eject_Signal_Debounce_0/ms_cnt[2]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74744, CLK => CLKINT_0_Y_0, Q
         => \Eject_Signal_Debounce_0/ms_cnt[2]_net_1\);
    
    \General_Controller_0/uc_send[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73768, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73601, Q => 
        \General_Controller_0_uc_send[1]\);
    
    HIEFFPLA_INST_0_67666 : AND3C
      port map(A => HIEFFPLA_NET_0_72843, B => 
        HIEFFPLA_NET_0_72816, C => HIEFFPLA_NET_0_72814, Y => 
        HIEFFPLA_NET_0_72829);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[2]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72801, Q => 
        \Sensors_0_acc_x[2]\);
    
    HIEFFPLA_INST_0_60128 : AO1D
      port map(A => HIEFFPLA_NET_0_74450, B => 
        HIEFFPLA_NET_0_74439, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74457);
    
    HIEFFPLA_INST_0_65011 : AO1B
      port map(A => HIEFFPLA_NET_0_73450, B => 
        HIEFFPLA_NET_0_73477, C => HIEFFPLA_NET_0_73482, Y => 
        HIEFFPLA_NET_0_73489);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/num_bytes_1[2]\ : 
        DFN1E1
      port map(D => HIEFFPLA_NET_0_72558, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72549, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_num_bytes[2]\);
    
    HIEFFPLA_INST_0_60081 : MX2
      port map(A => \Science_0_chan3_data[2]\, B => 
        \Science_0_chan3_data[6]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74464);
    
    HIEFFPLA_INST_0_70792 : NAND3C
      port map(A => HIEFFPLA_NET_0_72011, B => 
        HIEFFPLA_NET_0_72368, C => HIEFFPLA_NET_0_72371, Y => 
        HIEFFPLA_NET_0_72378);
    
    HIEFFPLA_INST_0_61669 : MX2
      port map(A => \SweepTable_0_RD[1]\, B => 
        \SweepTable_1_RD[1]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74163);
    
    HIEFFPLA_INST_0_61118 : AX1
      port map(A => HIEFFPLA_NET_0_74330, B => 
        HIEFFPLA_NET_0_74271, C => LED2_c, Y => 
        HIEFFPLA_NET_0_74272);
    
    \General_Controller_0/sweep_table_sweep_cnt[10]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74143, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[10]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72538, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/data_out[3]\ : 
        DFN0E1C1
      port map(D => ACCE_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73122, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\);
    
    \Communications_0/UART_0/tx_byte[3]\ : DFN1E1
      port map(D => \GS_Readout_0_send[3]\, CLK => CLKINT_0_Y_0, 
        E => HIEFFPLA_NET_0_75504, Q => 
        \Communications_0/UART_0/tx_byte[3]_net_1\);
    
    HIEFFPLA_INST_0_58828 : NOR3B
      port map(A => HIEFFPLA_NET_0_74645, B => 
        HIEFFPLA_NET_0_74432, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74678);
    
    \General_Controller_0/uc_tx_state[4]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73569, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[4]_net_1\);
    
    \CU_SYNC_pad/U0/U1\ : IOIN_IB
      port map(YIN => \CU_SYNC_pad/U0/NET1\, Y => CU_SYNC_c);
    
    \Science_0/ADC_READ_0/newflag\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73238, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73242, Q => 
        \Science_0/ADC_READ_0/newflag_net_1\);
    
    HIEFFPLA_INST_0_61897 : NOR3B
      port map(A => \General_Controller_0/uc_rx_byte[2]_net_1\, B
         => HIEFFPLA_NET_0_74082, C => 
        \General_Controller_0/uc_rx_byte[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74104);
    
    HIEFFPLA_INST_0_56921 : MX2
      port map(A => HIEFFPLA_NET_0_74984, B => 
        HIEFFPLA_NET_0_74912, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75195);
    
    HIEFFPLA_INST_0_57249 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[56]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_75114);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRYSYNC[3]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_14_Q\, 
        CLK => CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[3]\\\\\);
    
    HIEFFPLA_INST_0_68940 : NOR3A
      port map(A => HIEFFPLA_NET_0_72514, B => 
        HIEFFPLA_NET_0_72551, C => HIEFFPLA_NET_0_72501, Y => 
        HIEFFPLA_NET_0_72517);
    
    HIEFFPLA_INST_0_68368 : AND2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_i2c_repeat_start\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72668);
    
    HIEFFPLA_INST_0_62312 : AND3
      port map(A => HIEFFPLA_NET_0_73908, B => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, C => 
        HIEFFPLA_NET_0_73805, Y => HIEFFPLA_NET_0_74008);
    
    HIEFFPLA_INST_0_58473 : AOI1
      port map(A => HIEFFPLA_NET_0_74757, B => 
        HIEFFPLA_NET_0_74766, C => HIEFFPLA_NET_0_74756, Y => 
        HIEFFPLA_NET_0_74758);
    
    HIEFFPLA_INST_0_70767 : AOI1
      port map(A => HIEFFPLA_NET_0_72016, B => 
        HIEFFPLA_NET_0_72268, C => HIEFFPLA_NET_0_72234, Y => 
        HIEFFPLA_NET_0_72203);
    
    HIEFFPLA_INST_0_69913 : AND2B
      port map(A => HIEFFPLA_NET_0_72229, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72268);
    
    HIEFFPLA_INST_0_60532 : AND2A
      port map(A => \GS_Readout_0/subState[2]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74400);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[10]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72283, Q => 
        \Sensors_0_pressure_temp_raw[10]\);
    
    HIEFFPLA_INST_0_67955 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        B => HIEFFPLA_NET_0_72757, C => HIEFFPLA_NET_0_72775, Y
         => HIEFFPLA_NET_0_72767);
    
    \General_Controller_0/en_sensors\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74312, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => General_Controller_0_en_sensors);
    
    \General_Controller_0/uc_send[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73763, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73601, Q => 
        \General_Controller_0_uc_send[6]\);
    
    \General_Controller_0/status_bits_1[57]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74189, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[57]\);
    
    HIEFFPLA_INST_0_70556 : NOR3B
      port map(A => \Timing_0/m_count[6]_net_1\, B => 
        HIEFFPLA_NET_0_72084, C => \Timing_0/m_count[7]_net_1\, Y
         => HIEFFPLA_NET_0_72081);
    
    HIEFFPLA_INST_0_66990 : AOI1C
      port map(A => HIEFFPLA_NET_0_72980, B => 
        HIEFFPLA_NET_0_72978, C => HIEFFPLA_NET_0_72984, Y => 
        HIEFFPLA_NET_0_72989);
    
    \General_Controller_0/mission_mode\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74270, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/mission_mode_net_1\);
    
    HIEFFPLA_INST_0_55426 : AXOI4
      port map(A => HIEFFPLA_NET_0_75501, B => 
        \Communications_0/UART_0/tx_clk_count[0]_net_1\, C => 
        \Communications_0/UART_0/tx_clk_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75516);
    
    HIEFFPLA_INST_0_68101 : MX2B
      port map(A => HIEFFPLA_NET_0_72727, B => 
        HIEFFPLA_NET_0_72725, S => HIEFFPLA_NET_0_72878, Y => 
        HIEFFPLA_NET_0_72729);
    
    HIEFFPLA_INST_0_56046 : XNOR2
      port map(A => HIEFFPLA_NET_0_75279, B => 
        HIEFFPLA_NET_0_75294, Y => HIEFFPLA_NET_0_75360);
    
    HIEFFPLA_INST_0_60829 : XA1B
      port map(A => HIEFFPLA_NET_0_74347, B => 
        \GS_Readout_0/subState[4]_net_1\, C => 
        HIEFFPLA_NET_0_74350, Y => HIEFFPLA_NET_0_74351);
    
    HIEFFPLA_INST_0_59563 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[57]\, B => 
        \Data_Hub_Packets_0_status_packet[61]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74537);
    
    HIEFFPLA_INST_0_70710 : AND3
      port map(A => HIEFFPLA_NET_0_72034, B => 
        HIEFFPLA_NET_0_72033, C => \Timing_0/s_time[6]_net_1\, Y
         => HIEFFPLA_NET_0_72035);
    
    HIEFFPLA_INST_0_70605 : XOR2
      port map(A => \Timing_0/m_time[0]_net_1\, B => 
        HIEFFPLA_NET_0_72083, Y => HIEFFPLA_NET_0_72067);
    
    HIEFFPLA_INST_0_62947 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[3]_net_1\, 
        B => \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73860);
    
    \Science_0/ADC_READ_0/exp_packet_1[47]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[13]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[47]\);
    
    HIEFFPLA_INST_0_67242 : AND3
      port map(A => HIEFFPLA_NET_0_72749, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        C => HIEFFPLA_NET_0_72736, Y => HIEFFPLA_NET_0_72930);
    
    HIEFFPLA_INST_0_66740 : NOR2A
      port map(A => ACCE_SCL_c, B => 
        \Sensors_0/Accelerometer_0/state[8]\, Y => 
        HIEFFPLA_NET_0_73049);
    
    HIEFFPLA_INST_0_59481 : AO1D
      port map(A => HIEFFPLA_NET_0_74637, B => 
        \GS_Readout_0/subState[1]_net_1\, C => 
        HIEFFPLA_NET_0_74456, Y => HIEFFPLA_NET_0_74548);
    
    HIEFFPLA_INST_0_68369 : AND2
      port map(A => HIEFFPLA_NET_0_72700, B => 
        HIEFFPLA_NET_0_72698, Y => HIEFFPLA_NET_0_72667);
    
    HIEFFPLA_INST_0_70552 : NOR3B
      port map(A => \Timing_0/m_count[4]_net_1\, B => 
        HIEFFPLA_NET_0_72085, C => \Timing_0/m_count[1]_net_1\, Y
         => HIEFFPLA_NET_0_72082);
    
    HIEFFPLA_INST_0_62841 : AND3A
      port map(A => HIEFFPLA_NET_0_73810, B => 
        \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73885);
    
    HIEFFPLA_INST_0_56357 : AX1A
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, B
         => HIEFFPLA_NET_0_75350, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, Y
         => HIEFFPLA_NET_0_75302);
    
    HIEFFPLA_INST_0_64679 : AND2
      port map(A => 
        \General_Controller_0/uc_tx_nextstate[7]_net_1\, B => 
        HIEFFPLA_NET_0_73584, Y => HIEFFPLA_NET_0_73566);
    
    HIEFFPLA_INST_0_64463 : MX2A
      port map(A => \General_Controller_0/uc_tx_state[12]_net_1\, 
        B => HIEFFPLA_NET_0_73620, S => HIEFFPLA_NET_0_73561, Y
         => HIEFFPLA_NET_0_73621);
    
    HIEFFPLA_INST_0_64237 : MX2
      port map(A => HIEFFPLA_NET_0_73742, B => 
        HIEFFPLA_NET_0_73734, S => HIEFFPLA_NET_0_73588, Y => 
        HIEFFPLA_NET_0_73646);
    
    HIEFFPLA_INST_0_68675 : AO1
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[0]_net_1\, B
         => \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_72592);
    
    HIEFFPLA_INST_0_63242 : NOR3B
      port map(A => HIEFFPLA_NET_0_73780, B => 
        HIEFFPLA_NET_0_73907, C => HIEFFPLA_NET_0_73788, Y => 
        HIEFFPLA_NET_0_73800);
    
    HIEFFPLA_INST_0_55190 : AND3
      port map(A => \Communications_0/UART_0/rx_count[2]_net_1\, 
        B => \Communications_0/UART_0/rx_count[1]_net_1\, C => 
        \Communications_0/UART_0/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75564);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[7]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72800, Q => 
        \Sensors_0_acc_x[7]\);
    
    HIEFFPLA_INST_0_65788 : AO1A
      port map(A => \Science_0/ADC_READ_0/countere\, B => 
        HIEFFPLA_NET_0_73235, C => HIEFFPLA_NET_0_73280, Y => 
        HIEFFPLA_NET_0_73279);
    
    HIEFFPLA_INST_0_63106 : AND2
      port map(A => HIEFFPLA_NET_0_74026, B => 
        HIEFFPLA_NET_0_74070, Y => HIEFFPLA_NET_0_73827);
    
    HIEFFPLA_INST_0_68877 : AOI1
      port map(A => HIEFFPLA_NET_0_72527, B => 
        HIEFFPLA_NET_0_72486, C => HIEFFPLA_NET_0_72520, Y => 
        HIEFFPLA_NET_0_72534);
    
    HIEFFPLA_INST_0_71431 : OA1C
      port map(A => HIEFFPLA_NET_0_71968, B => 
        \Science_0/ADC_READ_0_G2[1]\, C => HIEFFPLA_NET_0_71995, 
        Y => HIEFFPLA_NET_0_73260);
    
    HIEFFPLA_INST_0_65404 : OR3B
      port map(A => \Science_0/ADC_READ_0/cnt2dn[5]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2dn[6]_net_1\, C => 
        HIEFFPLA_NET_0_73379, Y => HIEFFPLA_NET_0_73386);
    
    \General_Controller_0/uc_wen\ : DFN1E0C1
      port map(D => Communications_0_uc_tx_rdy, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73545, Q => General_Controller_0_uc_wen);
    
    HIEFFPLA_INST_0_55287 : AND2B
      port map(A => HIEFFPLA_NET_0_75583, B => 
        \Communications_0/UART_0/rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75545);
    
    HIEFFPLA_INST_0_64121 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_1[8]_net_1\, 
        B => 
        \General_Controller_0/constant_bias_voltage_1[0]_net_1\, 
        S => HIEFFPLA_NET_0_73558, Y => HIEFFPLA_NET_0_73665);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[5]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72464, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[5]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[2]\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72298, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72221, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[2]_net_1\);
    
    HIEFFPLA_INST_0_55656 : AND3
      port map(A => \Communications_0/UART_1/rx_count[2]_net_1\, 
        B => \Communications_0/UART_1/rx_count[1]_net_1\, C => 
        \Communications_0/UART_1/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75453);
    
    \Science_0/ADC_READ_0/exp_packet_1[34]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[0]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[34]\);
    
    HIEFFPLA_INST_0_61049 : NOR3B
      port map(A => HIEFFPLA_NET_0_74284, B => 
        \General_Controller_0/flight_state[4]_net_1\, C => 
        HIEFFPLA_NET_0_74281, Y => HIEFFPLA_NET_0_74287);
    
    HIEFFPLA_INST_0_64818 : AND3
      port map(A => HIEFFPLA_NET_0_73780, B => 
        HIEFFPLA_NET_0_74013, C => HIEFFPLA_NET_0_73533, Y => 
        HIEFFPLA_NET_0_73534);
    
    HIEFFPLA_INST_0_63220 : AND3
      port map(A => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, B => 
        HIEFFPLA_NET_0_74081, C => 
        \General_Controller_0/uc_rx_byte[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73803);
    
    HIEFFPLA_INST_0_58117 : AND2
      port map(A => \Science_0_exp_packet_0[37]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        Y => HIEFFPLA_NET_0_74847);
    
    HIEFFPLA_INST_0_57206 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[49]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75130);
    
    \Communications_0/UART_0/recv[1]\ : DFN1E1C1
      port map(D => \Communications_0/UART_0/rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75551, Q => 
        \Communications_0/UART_0_recv[1]\);
    
    HIEFFPLA_INST_0_55355 : AND3
      port map(A => \Communications_0/UART_0/tx_clk_count_i_0[5]\, 
        B => \Communications_0/UART_0/tx_clk_count_i_0[7]\, C => 
        \Communications_0/UART_0/tx_clk_count_i_0[6]\, Y => 
        HIEFFPLA_NET_0_75531);
    
    HIEFFPLA_INST_0_70795 : AOI1B
      port map(A => HIEFFPLA_NET_0_72540, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        C => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72010);
    
    HIEFFPLA_INST_0_57578 : AOI1
      port map(A => \Science_0_exp_packet_0[42]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74806, Y => HIEFFPLA_NET_0_75003);
    
    HIEFFPLA_INST_0_57667 : AO1
      port map(A => \Sensors_0_pressure_raw[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74790, Y => HIEFFPLA_NET_0_74976);
    
    HIEFFPLA_INST_0_57000 : AND3C
      port map(A => HIEFFPLA_NET_0_74867, B => 
        HIEFFPLA_NET_0_75046, C => HIEFFPLA_NET_0_74890, Y => 
        HIEFFPLA_NET_0_75184);
    
    HIEFFPLA_INST_0_55021 : XOR2
      port map(A => \General_Controller_0_unit_id[6]\, B => 
        \Communications_0/UART_0_recv[6]\, Y => 
        HIEFFPLA_NET_0_75613);
    
    \Science_0/SET_LP_GAIN_0/L2WR\ : DFN0C1
      port map(D => \Science_0/SET_LP_GAIN_0/state_i_0[2]\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => L2WR_c);
    
    HIEFFPLA_INST_0_71367 : OA1C
      port map(A => HIEFFPLA_NET_0_71969, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, C
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72004);
    
    HIEFFPLA_INST_0_70288 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        B => HIEFFPLA_NET_0_72180, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72181);
    
    HIEFFPLA_INST_0_69428 : MIN3X
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[2]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72391);
    
    HIEFFPLA_INST_0_57847 : AO1B
      port map(A => \Sensors_0_mag_time[20]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74926, Y => HIEFFPLA_NET_0_74927);
    
    HIEFFPLA_INST_0_60379 : MX2
      port map(A => \Science_0_chan4_data[4]\, B => 
        \Science_0_chan4_data[8]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74424);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[16]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[16]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[16]\);
    
    HIEFFPLA_INST_0_66219 : XO1
      port map(A => \Science_0/SET_LP_GAIN_0/old_G2[0]_net_1\, B
         => \Science_0/ADC_READ_0_G2[0]\, C => 
        HIEFFPLA_NET_0_73174, Y => HIEFFPLA_NET_0_73175);
    
    HIEFFPLA_INST_0_67752 : AO1A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        B => HIEFFPLA_NET_0_72736, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72809);
    
    \Science_0/ADC_READ_0/data_b[8]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[8]_net_1\);
    
    HIEFFPLA_INST_0_66309 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[2]\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73149);
    
    \General_Controller_0/sweep_table_sample_skip[9]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[9]_net_1\);
    
    HIEFFPLA_INST_0_70348 : AOI1D
      port map(A => General_Controller_0_st_ren1, B => 
        \SweepTable_0/WEBP\, C => 
        \General_Controller_0_st_raddr_1[6]\, Y => 
        \TableSelect_0_RADDR[6]\);
    
    HIEFFPLA_INST_0_64722 : OR3A
      port map(A => 
        \General_Controller_0/uc_tx_substate[0]_net_1\, B => 
        \General_Controller_0/uc_tx_substate[2]_net_1\, C => 
        HIEFFPLA_NET_0_73557, Y => HIEFFPLA_NET_0_73552);
    
    HIEFFPLA_INST_0_66042 : XA1B
      port map(A => HIEFFPLA_NET_0_73204, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, C => 
        \Science_0/DAC_SET_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73228);
    
    HIEFFPLA_INST_0_70361 : AND3
      port map(A => \Timekeeper_0_microseconds[19]\, B => 
        HIEFFPLA_NET_0_72158, C => 
        \Timekeeper_0_microseconds[20]\, Y => 
        HIEFFPLA_NET_0_72160);
    
    HIEFFPLA_INST_0_70132 : AO1
      port map(A => HIEFFPLA_NET_0_72192, B => 
        HIEFFPLA_NET_0_72181, C => HIEFFPLA_NET_0_72183, Y => 
        HIEFFPLA_NET_0_72212);
    
    HIEFFPLA_INST_0_64597 : NOR3A
      port map(A => HIEFFPLA_NET_0_73591, B => 
        HIEFFPLA_NET_0_73603, C => 
        \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73592);
    
    HIEFFPLA_INST_0_55416 : NAND2B
      port map(A => HIEFFPLA_NET_0_75517, B => 
        HIEFFPLA_NET_0_75527, Y => HIEFFPLA_NET_0_75518);
    
    HIEFFPLA_INST_0_65731 : NAND3
      port map(A => HIEFFPLA_NET_0_73295, B => 
        \Science_0/ADC_READ_0/cnt_chan[0]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt_chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73296);
    
    HIEFFPLA_INST_0_62875 : AO1A
      port map(A => HIEFFPLA_NET_0_74071, B => 
        HIEFFPLA_NET_0_73956, C => HIEFFPLA_NET_0_73876, Y => 
        HIEFFPLA_NET_0_73877);
    
    \TOP_UART_RX_pad/U0/U0\ : IOPAD_IN
      port map(PAD => TOP_UART_RX, Y => \TOP_UART_RX_pad/U0/NET1\);
    
    HIEFFPLA_INST_0_57254 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[61]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_75109);
    
    HIEFFPLA_INST_0_70476 : AND3
      port map(A => \Timekeeper_0_milliseconds[13]\, B => 
        HIEFFPLA_NET_0_72127, C => 
        \Timekeeper_0_milliseconds[14]\, Y => 
        HIEFFPLA_NET_0_72118);
    
    HIEFFPLA_INST_0_69477 : OR3A
      port map(A => PRESSURE_SCL_c, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        C => HIEFFPLA_NET_0_72344, Y => HIEFFPLA_NET_0_72379);
    
    \Science_0/ADC_READ_0/cnt1up[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73392, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1up[3]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/data_out[26]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75217, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[26]\);
    
    HIEFFPLA_INST_0_67428 : NAND3C
      port map(A => HIEFFPLA_NET_0_72791, B => 
        HIEFFPLA_NET_0_72743, C => HIEFFPLA_NET_0_72891, Y => 
        HIEFFPLA_NET_0_72883);
    
    HIEFFPLA_INST_0_60165 : MX2
      port map(A => \Sensors_0_pressure_raw[19]\, B => 
        \Sensors_0_pressure_raw[23]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74451);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[0]\ : 
        DFN0E1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        CLK => ClockDivs_0_clk_800kHz, E => HIEFFPLA_NET_0_72354, 
        Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[0]_net_1\);
    
    HIEFFPLA_INST_0_69395 : NOR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => HIEFFPLA_NET_0_72351, C => HIEFFPLA_NET_0_72423, Y
         => HIEFFPLA_NET_0_72399);
    
    \General_Controller_0/gs_id[3]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73922, Q => 
        \General_Controller_0_gs_id[3]\);
    
    HIEFFPLA_INST_0_88369 : AO18
      port map(A => HIEFFPLA_NET_0_75321, B => 
        HIEFFPLA_NET_0_75320, C => HIEFFPLA_NET_0_75304, Y => 
        HIEFFPLA_NET_0_88384);
    
    HIEFFPLA_INST_0_65758 : AND2A
      port map(A => HIEFFPLA_NET_0_73241, B => 
        HIEFFPLA_NET_0_73286, Y => HIEFFPLA_NET_0_73287);
    
    HIEFFPLA_INST_0_55683 : XNOR2
      port map(A => \Communications_0/UART_1/rx_count[1]_net_1\, 
        B => \Communications_0/UART_1/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75447);
    
    HIEFFPLA_INST_0_61113 : AX1
      port map(A => HIEFFPLA_NET_0_74334, B => 
        HIEFFPLA_NET_0_74326, C => LED1_c, Y => 
        HIEFFPLA_NET_0_74273);
    
    HIEFFPLA_INST_0_55799 : MX2C
      port map(A => \Communications_0/UART_1/tx_byte[0]_net_1\, B
         => \Communications_0/UART_1/tx_byte[4]_net_1\, S => 
        \Communications_0/UART_1/tx_count[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75424);
    
    AFLSDF_INV_30 : INV
      port map(A => General_Controller_0_status_new_data, Y => 
        \AFLSDF_INV_30\);
    
    HIEFFPLA_INST_0_55709 : AOI1D
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\, B => 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\, C => 
        HIEFFPLA_NET_0_75444, Y => HIEFFPLA_NET_0_75440);
    
    HIEFFPLA_INST_0_67364 : NAND3C
      port map(A => HIEFFPLA_NET_0_72933, B => 
        HIEFFPLA_NET_0_72892, C => HIEFFPLA_NET_0_72927, Y => 
        HIEFFPLA_NET_0_72897);
    
    HIEFFPLA_INST_0_55306 : MX2
      port map(A => HIEFFPLA_NET_0_75540, B => 
        HIEFFPLA_NET_0_75539, S => 
        \Communications_0/UART_0/tx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75542);
    
    \LED2_pad/U0/U0\ : IOPAD_TRI
      port map(D => \LED2_pad/U0/NET1\, E => \LED2_pad/U0/NET2\, 
        PAD => LED2);
    
    HIEFFPLA_INST_0_55922 : NOR3B
      port map(A => \Communications_0/UART_1/tx_state[1]_net_1\, 
        B => \Communications_0/UART_1/tx_count[2]_net_1\, C => 
        \Communications_0/UART_1/tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75394);
    
    \Data_Saving_0/Packet_Saver_0/data_out[2]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75213, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[2]\);
    
    HIEFFPLA_INST_0_58397 : AO1
      port map(A => \Sensors_0_mag_x[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_75098, Y => HIEFFPLA_NET_0_74780);
    
    HIEFFPLA_INST_0_70491 : XOR2
      port map(A => HIEFFPLA_NET_0_72127, B => 
        \Timekeeper_0_milliseconds[13]\, Y => 
        HIEFFPLA_NET_0_72112);
    
    HIEFFPLA_INST_0_67239 : AOI1C
      port map(A => HIEFFPLA_NET_0_72904, B => 
        HIEFFPLA_NET_0_72899, C => HIEFFPLA_NET_0_72902, Y => 
        HIEFFPLA_NET_0_72931);
    
    \Communications_0/UART_1/recv[3]\ : DFN1E1C1
      port map(D => \Communications_0/UART_1/rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75441, Q => \Communications_0_uc_recv[3]\);
    
    \General_Controller_0/constant_bias_voltage_1[1]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[1]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[1]_net_1\);
    
    HIEFFPLA_INST_0_64882 : AND3B
      port map(A => \I2C_PassThrough_0/cnt[0]_net_1\, B => 
        \I2C_PassThrough_0/cnt[3]_net_1\, C => 
        HIEFFPLA_NET_0_73519, Y => HIEFFPLA_NET_0_73518);
    
    \General_Controller_0/constant_bias_voltage_0[10]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[10]_net_1\);
    
    \Science_0/ADC_READ_0/cnt4dn[2]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73316, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4dn[2]_net_1\);
    
    HIEFFPLA_INST_0_57248 : AND2
      port map(A => \Sensors_0_acc_time[15]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, Y
         => HIEFFPLA_NET_0_75115);
    
    HIEFFPLA_INST_0_68892 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        Y => HIEFFPLA_NET_0_72530);
    
    HIEFFPLA_INST_0_57475 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_75034, Y => HIEFFPLA_NET_0_75035);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[9]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72753, Q => 
        \Sensors_0_acc_z[9]\);
    
    HIEFFPLA_INST_0_65695 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt4up[2]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt4up[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt4up[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73307);
    
    \Science_0/ADC_READ_0/chan4_data[10]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[10]\);
    
    \Data_Saving_0/Packet_Saver_0/data_out[20]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75224, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[20]\);
    
    HIEFFPLA_INST_0_70680 : AX1C
      port map(A => HIEFFPLA_NET_0_72034, B => 
        HIEFFPLA_NET_0_72033, C => \Timing_0/s_time[4]_net_1\, Y
         => HIEFFPLA_NET_0_72046);
    
    HIEFFPLA_INST_0_58572 : AX1
      port map(A => HIEFFPLA_NET_0_74739, B => 
        HIEFFPLA_NET_0_74737, C => 
        \Eject_Signal_Debounce_0/ms_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74732);
    
    HIEFFPLA_INST_0_57286 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[46]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75094);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1E1C0_data_out[3]\\\\/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75284, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \FMC_DA_c[3]\);
    
    HIEFFPLA_INST_0_68549 : NAND2B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[5]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72620);
    
    HIEFFPLA_INST_0_59854 : MX2
      port map(A => \ch3_data_net_0[8]\, B => 
        \Sensors_0_acc_z[0]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74497);
    
    HIEFFPLA_INST_0_58980 : NOR3B
      port map(A => HIEFFPLA_NET_0_74617, B => 
        HIEFFPLA_NET_0_74394, C => HIEFFPLA_NET_0_74397, Y => 
        HIEFFPLA_NET_0_74644);
    
    HIEFFPLA_INST_0_70180 : NOR3B
      port map(A => HIEFFPLA_NET_0_72285, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        C => HIEFFPLA_NET_0_72284, Y => HIEFFPLA_NET_0_72200);
    
    \Sensors_0/Gyro_0/I2C_Master_0/state[0]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72615, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\);
    
    \LA1_pad/U0/U0\ : IOPAD_TRI
      port map(D => \LA1_pad/U0/NET1\, E => \LA1_pad/U0/NET2\, 
        PAD => LA1);
    
    \Science_0/ADC_READ_0/chan5_data[7]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[7]\);
    
    \ClockDivs_0/cnt_800kHz[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75628, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \ClockDivs_0/cnt_800kHz[3]_net_1\);
    
    \General_Controller_0/sweep_table_samples_per_point[0]\ : 
        DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[0]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[0]_net_1\);
    
    HIEFFPLA_INST_0_66458 : AND3A
      port map(A => HIEFFPLA_NET_0_73143, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        C => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73115);
    
    HIEFFPLA_INST_0_60629 : MX2
      port map(A => \Science_0_chan0_data[7]\, B => 
        \Science_0_chan0_data[11]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74384);
    
    HIEFFPLA_INST_0_61155 : OR3A
      port map(A => \General_Controller_0/state_seconds[7]_net_1\, 
        B => HIEFFPLA_NET_0_74248, C => HIEFFPLA_NET_0_74245, Y
         => HIEFFPLA_NET_0_74261);
    
    HIEFFPLA_INST_0_56742 : MX2B
      port map(A => HIEFFPLA_NET_0_75184, B => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[1]_net_1\, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75218);
    
    HIEFFPLA_INST_0_66174 : MX2B
      port map(A => \Science_0/DAC_SET_0/vector[7]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73188);
    
    HIEFFPLA_INST_0_66094 : AND3C
      port map(A => HIEFFPLA_NET_0_73208, B => 
        HIEFFPLA_NET_0_73231, C => HIEFFPLA_NET_0_73211, Y => 
        HIEFFPLA_NET_0_73210);
    
    HIEFFPLA_INST_0_57740 : AOI1
      port map(A => \Science_0_exp_packet_0[60]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74818, Y => HIEFFPLA_NET_0_74956);
    
    HIEFFPLA_INST_0_57090 : AOI1
      port map(A => \Sensors_0_pressure_raw[22]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, C
         => HIEFFPLA_NET_0_74884, Y => HIEFFPLA_NET_0_75169);
    
    HIEFFPLA_INST_0_55653 : NOR2A
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[28]_net_1\, B => 
        HIEFFPLA_NET_0_75467, Y => HIEFFPLA_NET_0_75454);
    
    \General_Controller_0/uc_rx_byte[7]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[7]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte[7]_net_1\);
    
    HIEFFPLA_INST_0_67297 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72914);
    
    HIEFFPLA_INST_0_55527 : AND2B
      port map(A => \Communications_0/UART_1/rx_count[2]_net_1\, 
        B => \Communications_0/UART_1/rx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75487);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[14]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[14]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[14]\);
    
    HIEFFPLA_INST_0_66889 : AND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73010);
    
    HIEFFPLA_INST_0_57343 : AOI1
      port map(A => \Science_0_exp_packet_0[12]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_75070, Y => HIEFFPLA_NET_0_75071);
    
    HIEFFPLA_INST_0_69473 : AOI1
      port map(A => HIEFFPLA_NET_0_72355, B => PRESSURE_SCL_c, C
         => HIEFFPLA_NET_0_72342, Y => HIEFFPLA_NET_0_72380);
    
    \Sensors_0/Gyro_0/I2C_Master_0/s_ack_error\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72630, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72665, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_s_ack_error\);
    
    \Science_0/DAC_SET_0/CS\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_73227, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => LDCS_c);
    
    HIEFFPLA_INST_0_65234 : OR3B
      port map(A => \Sensors_0_pressure_raw[22]\, B => 
        \Sensors_0_pressure_raw[20]\, C => HIEFFPLA_NET_0_73440, 
        Y => HIEFFPLA_NET_0_73438);
    
    HIEFFPLA_INST_0_60747 : MX2
      port map(A => \Science_0_chan5_data[11]\, B => 
        \Science_0_chan4_data[3]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74364);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[4]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[4]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[4]\);
    
    HIEFFPLA_INST_0_66390 : NAND3C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73131);
    
    HIEFFPLA_INST_0_64197 : AOI1C
      port map(A => \General_Controller_0/uc_tx_state[14]_net_1\, 
        B => HIEFFPLA_NET_0_73747, C => 
        \General_Controller_0/uc_tx_state[12]_net_1\, Y => 
        HIEFFPLA_NET_0_73651);
    
    HIEFFPLA_INST_0_67631 : AOI1C
      port map(A => HIEFFPLA_NET_0_72894, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        C => HIEFFPLA_NET_0_72837, Y => HIEFFPLA_NET_0_72838);
    
    HIEFFPLA_INST_0_65947 : OA1C
      port map(A => HIEFFPLA_NET_0_73252, B => 
        \Science_0/ADC_READ_0_G3[1]\, C => HIEFFPLA_NET_0_73350, 
        Y => HIEFFPLA_NET_0_73254);
    
    HIEFFPLA_INST_0_68852 : NAND3C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, B
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, Y
         => HIEFFPLA_NET_0_72540);
    
    HIEFFPLA_INST_0_59002 : NOR3B
      port map(A => HIEFFPLA_NET_0_74615, B => 
        HIEFFPLA_NET_0_74436, C => HIEFFPLA_NET_0_74510, Y => 
        HIEFFPLA_NET_0_74639);
    
    HIEFFPLA_INST_0_58508 : NAND2B
      port map(A => HIEFFPLA_NET_0_74745, B => 
        HIEFFPLA_NET_0_74740, Y => HIEFFPLA_NET_0_74746);
    
    HIEFFPLA_INST_0_55912 : NOR3A
      port map(A => 
        \Communications_0/UART_1/tx_clk_count[1]_net_1\, B => 
        \Communications_0/UART_1/tx_state[0]_net_1\, C => 
        \Communications_0/UART_1/tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75397);
    
    \FPGA_BUF_INT_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => FPGA_BUF_INT_c, E => \VCC\, DOUT => 
        \FPGA_BUF_INT_pad/U0/NET1\, EOUT => 
        \FPGA_BUF_INT_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_56976 : MX2
      port map(A => HIEFFPLA_NET_0_74964, B => 
        HIEFFPLA_NET_0_74894, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75188);
    
    \Communications_0/UART_1/tx_count[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75391, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75388, Q => 
        \Communications_0/UART_1/tx_count[2]_net_1\);
    
    HIEFFPLA_INST_0_60146 : MX2
      port map(A => HIEFFPLA_NET_0_74342, B => 
        HIEFFPLA_NET_0_74376, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74454);
    
    HIEFFPLA_INST_0_55270 : AND2B
      port map(A => HIEFFPLA_NET_0_75551, B => 
        HIEFFPLA_NET_0_75594, Y => HIEFFPLA_NET_0_75548);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[8]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72800, Q => 
        \Sensors_0_acc_x[8]\);
    
    HIEFFPLA_INST_0_61364 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[3]\, B => 
        UC_PWR_EN_c, S => HIEFFPLA_NET_0_74266, Y => 
        HIEFFPLA_NET_0_74208);
    
    HIEFFPLA_INST_0_55740 : MX2A
      port map(A => HIEFFPLA_NET_0_75378, B => 
        HIEFFPLA_NET_0_75482, S => 
        \Communications_0/UART_1/rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75434);
    
    HIEFFPLA_INST_0_55069 : AND3
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[25]_net_1\, B => 
        HIEFFPLA_NET_0_75586, C => 
        \Communications_0/UART_0/rx_clk_count[26]_net_1\, Y => 
        HIEFFPLA_NET_0_75598);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72461, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\);
    
    HIEFFPLA_INST_0_70458 : AND3
      port map(A => \Timekeeper_0_milliseconds[17]\, B => 
        HIEFFPLA_NET_0_72121, C => 
        \Timekeeper_0_milliseconds[18]\, Y => 
        HIEFFPLA_NET_0_72123);
    
    HIEFFPLA_INST_0_67040 : AOI1C
      port map(A => \Sensors_0/Accelerometer_0/state_0[8]\, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[1]\, 
        C => HIEFFPLA_NET_0_72890, Y => HIEFFPLA_NET_0_72981);
    
    HIEFFPLA_INST_0_57558 : AND2
      port map(A => \Sensors_0_gyro_time[20]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75009);
    
    HIEFFPLA_INST_0_56243 : XNOR3
      port map(A => HIEFFPLA_NET_0_75277, B => 
        HIEFFPLA_NET_0_75290, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\, Y
         => HIEFFPLA_NET_0_75326);
    
    HIEFFPLA_INST_0_57196 : AO1
      port map(A => \Sensors_0_pressure_time[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75092, Y => HIEFFPLA_NET_0_75133);
    
    HIEFFPLA_INST_0_66451 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => HIEFFPLA_NET_0_73116, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73117);
    
    HIEFFPLA_INST_0_59802 : AO1
      port map(A => HIEFFPLA_NET_0_74404, B => 
        HIEFFPLA_NET_0_74341, C => HIEFFPLA_NET_0_74505, Y => 
        HIEFFPLA_NET_0_74506);
    
    \Communications_0/UART_1/rx_clk_count[31]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75456, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75443, Q => 
        \Communications_0/UART_1/rx_clk_count_c0\);
    
    \General_Controller_0/uc_tx_substate[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73550, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_tx_substate[1]_net_1\);
    
    HIEFFPLA_INST_0_70031 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72242);
    
    HIEFFPLA_INST_0_64163 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_1[6]_net_1\, 
        B => 
        \General_Controller_0/constant_bias_voltage_1[14]_net_1\, 
        S => \General_Controller_0/uc_tx_substate[1]_net_1\, Y
         => HIEFFPLA_NET_0_73659);
    
    HIEFFPLA_INST_0_61323 : AND2B
      port map(A => HIEFFPLA_NET_0_74295, B => 
        HIEFFPLA_NET_0_74293, Y => HIEFFPLA_NET_0_74217);
    
    HIEFFPLA_INST_0_56072 : XA1
      port map(A => HIEFFPLA_NET_0_75259, B => 
        HIEFFPLA_NET_0_75323, C => HIEFFPLA_NET_0_75354, Y => 
        HIEFFPLA_NET_0_75355);
    
    \General_Controller_0/status_bits_1[42]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74204, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[42]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[22]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[22]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[22]\);
    
    HIEFFPLA_INST_0_57291 : AND2
      port map(A => \Sensors_0_gyro_time[12]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75089);
    
    HIEFFPLA_INST_0_55833 : NAND2
      port map(A => 
        \Communications_0/UART_1/tx_clk_count[1]_net_1\, B => 
        \Communications_0/UART_1/tx_clk_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75417);
    
    HIEFFPLA_INST_0_55592 : NOR3B
      port map(A => HIEFFPLA_NET_0_75476, B => 
        \Communications_0/UART_1/rx_clk_count[28]_net_1\, C => 
        \Communications_0/UART_1/rx_clk_count[27]_net_1\, Y => 
        HIEFFPLA_NET_0_75472);
    
    HIEFFPLA_INST_0_55506 : NOR3B
      port map(A => HIEFFPLA_NET_0_75485, B => 
        HIEFFPLA_NET_0_75488, C => 
        \Communications_0/UART_1/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75494);
    
    \Data_Saving_0/Packet_Saver_0/data_out[9]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75204, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[9]\);
    
    AFLSDF_INV_18 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_18\);
    
    HIEFFPLA_INST_0_69345 : AOI1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72413);
    
    HIEFFPLA_INST_0_60251 : OR3B
      port map(A => \GS_Readout_0/subState[4]_net_1\, B => 
        HIEFFPLA_NET_0_74636, C => HIEFFPLA_NET_0_74374, Y => 
        HIEFFPLA_NET_0_74441);
    
    HIEFFPLA_INST_0_55108 : AND2B
      port map(A => \Communications_0/UART_0/rx_state[1]_net_1\, 
        B => \Communications_0/UART_0/rx_clk_count[24]_net_1\, Y
         => HIEFFPLA_NET_0_75588);
    
    \FMC_DA_pad[0]/U0/U0\ : IOPAD_TRI
      port map(D => \FMC_DA_pad[0]/U0/NET1\, E => 
        \FMC_DA_pad[0]/U0/NET2\, PAD => FMC_DA(0));
    
    HIEFFPLA_INST_0_66330 : NOR3A
      port map(A => HIEFFPLA_NET_0_73148, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[3]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73144);
    
    HIEFFPLA_INST_0_64580 : OR3A
      port map(A => HIEFFPLA_NET_0_73592, B => 
        \General_Controller_0/uc_tx_state[0]_net_1\, C => 
        \General_Controller_0/uc_tx_state[14]_net_1\, Y => 
        HIEFFPLA_NET_0_73597);
    
    HIEFFPLA_INST_0_62623 : NAND3C
      port map(A => HIEFFPLA_NET_0_73941, B => 
        HIEFFPLA_NET_0_74037, C => HIEFFPLA_NET_0_74009, Y => 
        HIEFFPLA_NET_0_73942);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[9]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[9]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[9]\);
    
    HIEFFPLA_INST_0_70003 : AO1
      port map(A => HIEFFPLA_NET_0_72245, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        C => HIEFFPLA_NET_0_72247, Y => HIEFFPLA_NET_0_72249);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRYSYNC[7]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_13_Q\, 
        CLK => CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[7]\\\\\);
    
    HIEFFPLA_INST_0_64488 : NOR3A
      port map(A => \General_Controller_0/uc_tx_state[14]_net_1\, 
        B => Communications_0_uc_tx_rdy, C => 
        HIEFFPLA_NET_0_73558, Y => HIEFFPLA_NET_0_73616);
    
    \Communications_0/UART_1/tx_byte[0]\ : DFN1E1
      port map(D => \General_Controller_0_uc_send[0]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_75385, Q => 
        \Communications_0/UART_1/tx_byte[0]_net_1\);
    
    HIEFFPLA_INST_0_65047 : OA1C
      port map(A => \Sensors_0_pressure_raw[22]\, B => 
        HIEFFPLA_NET_0_73455, C => \Sensors_0_pressure_raw[23]\, 
        Y => HIEFFPLA_NET_0_73481);
    
    HIEFFPLA_INST_0_63426 : MX2
      port map(A => HIEFFPLA_NET_0_73756, B => 
        HIEFFPLA_NET_0_73690, S => HIEFFPLA_NET_0_73608, Y => 
        HIEFFPLA_NET_0_73764);
    
    HIEFFPLA_INST_0_69178 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, B
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        Y => HIEFFPLA_NET_0_72454);
    
    \LED1_pad/U0/U0\ : IOPAD_TRI
      port map(D => \LED1_pad/U0/NET1\, E => \LED1_pad/U0/NET2\, 
        PAD => LED1);
    
    HIEFFPLA_INST_0_68498 : AO1C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\, B => 
        HIEFFPLA_NET_0_72702, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_72636);
    
    HIEFFPLA_INST_0_62015 : XO1
      port map(A => 
        \General_Controller_0/uc_rx_prev_state[1]_net_1\, B => 
        \General_Controller_0/uc_rx_prev_state[2]_net_1\, C => 
        Communications_0_uc_rx_rdy, Y => HIEFFPLA_NET_0_74072);
    
    HIEFFPLA_INST_0_70879 : AX1D
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[0]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[1]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72007);
    
    HIEFFPLA_INST_0_66236 : XO1
      port map(A => \Science_0/SET_LP_GAIN_0/old_G3[1]_net_1\, B
         => \Science_0/ADC_READ_0_G3[1]\, C => 
        HIEFFPLA_NET_0_73170, Y => HIEFFPLA_NET_0_73171);
    
    HIEFFPLA_INST_0_60223 : MX2
      port map(A => HIEFFPLA_NET_0_74434, B => 
        HIEFFPLA_NET_0_74553, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74444);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_new_data\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72564, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, Q
         => Sensors_0_gyro_new_data);
    
    HIEFFPLA_INST_0_69126 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[5]_net_1\, 
        C => HIEFFPLA_NET_0_72556, Y => HIEFFPLA_NET_0_72465);
    
    \Communications_0/UART_0/tx_byte[4]\ : DFN1E1
      port map(D => \GS_Readout_0_send[4]\, CLK => CLKINT_0_Y_0, 
        E => HIEFFPLA_NET_0_75504, Q => 
        \Communications_0/UART_0/tx_byte[4]_net_1\);
    
    HIEFFPLA_INST_0_66664 : OR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        B => HIEFFPLA_NET_0_73070, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_73071);
    
    HIEFFPLA_INST_0_61213 : OR3B
      port map(A => \General_Controller_0/state_seconds[3]_net_1\, 
        B => \General_Controller_0/state_seconds[4]_net_1\, C => 
        HIEFFPLA_NET_0_74262, Y => HIEFFPLA_NET_0_74248);
    
    HIEFFPLA_INST_0_58285 : AO1
      port map(A => \Sensors_0_mag_x[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_75100, Y => HIEFFPLA_NET_0_74812);
    
    HIEFFPLA_INST_0_55640 : XA1A
      port map(A => HIEFFPLA_NET_0_75475, B => 
        \Communications_0/UART_1/rx_clk_count[29]_net_1\, C => 
        HIEFFPLA_NET_0_75437, Y => HIEFFPLA_NET_0_75458);
    
    \Timekeeper_0/microseconds[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72140, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[1]\);
    
    HIEFFPLA_INST_0_61931 : NAND3B
      port map(A => HIEFFPLA_NET_0_74016, B => 
        HIEFFPLA_NET_0_73808, C => HIEFFPLA_NET_0_74095, Y => 
        HIEFFPLA_NET_0_74096);
    
    HIEFFPLA_INST_0_64347 : MX2
      port map(A => HIEFFPLA_NET_0_73723, B => 
        HIEFFPLA_NET_0_73715, S => HIEFFPLA_NET_0_73619, Y => 
        HIEFFPLA_NET_0_73635);
    
    HIEFFPLA_INST_0_60731 : XA1
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, C => 
        HIEFFPLA_NET_0_74559, Y => HIEFFPLA_NET_0_74367);
    
    \Science_0/ADC_READ_0/cnt3up[1]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73335, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3up[1]_net_1\);
    
    HIEFFPLA_INST_0_70084 : OR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72225);
    
    HIEFFPLA_INST_0_59397 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[0]\, B => 
        \Data_Hub_Packets_0_status_packet[4]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74560);
    
    HIEFFPLA_INST_0_64958 : AND3
      port map(A => HIEFFPLA_NET_0_73501, B => 
        \I2C_PassThrough_0/cnt[2]_net_1\, C => 
        \I2C_PassThrough_0/cnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73503);
    
    \General_Controller_0/uc_rx_state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73997, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_state[1]_net_1\);
    
    HIEFFPLA_INST_0_67126 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[4]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72960);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[3]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72783, Q => 
        \Sensors_0_mag_y[3]\);
    
    HIEFFPLA_INST_0_61978 : NAND2
      port map(A => \General_Controller_0/uc_rx_byte[0]_net_1\, B
         => \General_Controller_0/uc_rx_byte[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74084);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[2]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72767, Q => 
        \Sensors_0_acc_y[2]\);
    
    HIEFFPLA_INST_0_61031 : AO1
      port map(A => HIEFFPLA_NET_0_74257, B => 
        \General_Controller_0/flight_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_74286, Y => HIEFFPLA_NET_0_74291);
    
    HIEFFPLA_INST_0_65511 : AND2
      port map(A => HIEFFPLA_NET_0_73351, B => 
        \Science_0/ADC_READ_0/cnt3dn[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73358);
    
    HIEFFPLA_INST_0_57310 : AND2
      port map(A => \Sensors_0_gyro_time[23]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75081);
    
    HIEFFPLA_INST_0_60581 : MX2A
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        HIEFFPLA_NET_0_74562, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74392);
    
    HIEFFPLA_INST_0_70806 : OA1A
      port map(A => HIEFFPLA_NET_0_72505, B => 
        HIEFFPLA_NET_0_72506, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, Y
         => HIEFFPLA_NET_0_72009);
    
    HIEFFPLA_INST_0_63370 : XA1
      port map(A => 
        \General_Controller_0/uc_rx_substate[4]_net_1\, B => 
        HIEFFPLA_NET_0_73534, C => HIEFFPLA_NET_0_73965, Y => 
        HIEFFPLA_NET_0_73770);
    
    HIEFFPLA_INST_0_58671 : NOR3A
      port map(A => HIEFFPLA_NET_0_74682, B => 
        HIEFFPLA_NET_0_74659, C => HIEFFPLA_NET_0_74626, Y => 
        HIEFFPLA_NET_0_74707);
    
    HIEFFPLA_INST_0_64669 : AND2
      port map(A => 
        \General_Controller_0/uc_tx_nextstate[2]_net_1\, B => 
        HIEFFPLA_NET_0_73584, Y => HIEFFPLA_NET_0_73571);
    
    HIEFFPLA_INST_0_69879 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        B => HIEFFPLA_NET_0_72239, C => HIEFFPLA_NET_0_72227, Y
         => HIEFFPLA_NET_0_72281);
    
    \Timekeeper_0/microseconds[9]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72128, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[9]\);
    
    HIEFFPLA_INST_0_62421 : NOR3A
      port map(A => HIEFFPLA_NET_0_74026, B => 
        HIEFFPLA_NET_0_73811, C => HIEFFPLA_NET_0_73804, Y => 
        HIEFFPLA_NET_0_73985);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_new_data\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73008, Q => Sensors_0_acc_new_data);
    
    HIEFFPLA_INST_0_70505 : XOR2
      port map(A => \Timekeeper_0_milliseconds[0]\, B => 
        \Timekeeper_0_milliseconds[1]\, Y => HIEFFPLA_NET_0_72105);
    
    HIEFFPLA_INST_0_67502 : AO1B
      port map(A => HIEFFPLA_NET_0_72778, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        C => HIEFFPLA_NET_0_72863, Y => HIEFFPLA_NET_0_72864);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[23]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[23]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[23]\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73138, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\);
    
    \Timekeeper_0/microseconds[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72135, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[2]\);
    
    HIEFFPLA_INST_0_63516 : MX2
      port map(A => HIEFFPLA_NET_0_73680, B => 
        HIEFFPLA_NET_0_73672, S => HIEFFPLA_NET_0_73621, Y => 
        HIEFFPLA_NET_0_73755);
    
    HIEFFPLA_INST_0_66758 : NAND2
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        B => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73043);
    
    HIEFFPLA_INST_0_59525 : MX2
      port map(A => HIEFFPLA_NET_0_74550, B => 
        HIEFFPLA_NET_0_74538, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74542);
    
    \SCIENCE_TX_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => SCIENCE_TX_c_c, E => \VCC\, DOUT => 
        \SCIENCE_TX_pad/U0/NET1\, EOUT => 
        \SCIENCE_TX_pad/U0/NET2\);
    
    \Science_0/ADC_READ_0/exp_packet_1[21]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[5]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[21]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/data_out_1[2]\ : 
        DFN1E1
      port map(D => HIEFFPLA_NET_0_73006, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72795, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[2]\);
    
    HIEFFPLA_INST_0_64481 : AND3B
      port map(A => 
        \General_Controller_0/constant_bias_probe_id[0]_net_1\, B
         => \General_Controller_0/un10_uc_tx_rdy_i[1]\, C => 
        \General_Controller_0/uc_tx_state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73618);
    
    \Communications_0/FFU_Command_Checker_0/command_out[5]\ : 
        DFN1E1C1
      port map(D => \Communications_0/UART_0_recv[5]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75625, Q => \Communications_0_ext_recv[5]\);
    
    HIEFFPLA_INST_0_68225 : MX2
      port map(A => HIEFFPLA_NET_0_72706, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_i2c_addr[0]\, S => 
        HIEFFPLA_NET_0_72702, Y => HIEFFPLA_NET_0_72700);
    
    HIEFFPLA_INST_0_68491 : OA1C
      port map(A => HIEFFPLA_NET_0_72620, B => 
        HIEFFPLA_NET_0_72705, C => HIEFFPLA_NET_0_72637, Y => 
        HIEFFPLA_NET_0_72638);
    
    \Science_0/ADC_READ_0/chan2_data[8]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[8]\);
    
    HIEFFPLA_INST_0_68458 : MX2
      port map(A => HIEFFPLA_NET_0_72657, B => 
        HIEFFPLA_NET_0_72656, S => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_72646);
    
    HIEFFPLA_INST_0_70766 : OR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72017);
    
    HIEFFPLA_INST_0_59933 : MX2
      port map(A => HIEFFPLA_NET_0_74483, B => 
        HIEFFPLA_NET_0_74545, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74486);
    
    HIEFFPLA_INST_0_60993 : AXOI5
      port map(A => \General_Controller_0/ext_rx_state_i_0[1]\, B
         => Communications_0_ext_rx_rdy, C => 
        \General_Controller_0/ext_rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74302);
    
    HIEFFPLA_INST_0_56531 : XOR2
      port map(A => HIEFFPLA_NET_0_75256, B => 
        \Data_Saving_0/Interrupt_Generator_0/counter[3]_net_1\, Y
         => HIEFFPLA_NET_0_75250);
    
    AFLSDF_INV_3 : INV
      port map(A => \Data_Saving_0/FPGA_Buffer_0/MEMRENEG\, Y => 
        \AFLSDF_INV_3\);
    
    \General_Controller_0/temp_first_byte[5]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73872, Q => 
        \General_Controller_0/temp_first_byte[5]_net_1\);
    
    HIEFFPLA_INST_0_66202 : XO1
      port map(A => \Science_0/SET_LP_GAIN_0/old_G1[1]_net_1\, B
         => \Science_0/ADC_READ_0_G1[1]\, C => 
        HIEFFPLA_NET_0_73178, Y => HIEFFPLA_NET_0_73179);
    
    HIEFFPLA_INST_0_66689 : AND3C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_73063);
    
    HIEFFPLA_INST_0_66413 : MX2
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[1]\, 
        S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_73126);
    
    HIEFFPLA_INST_0_68653 : AO1
      port map(A => HIEFFPLA_NET_0_72590, B => 
        HIEFFPLA_NET_0_72669, C => HIEFFPLA_NET_0_72587, Y => 
        HIEFFPLA_NET_0_72596);
    
    HIEFFPLA_INST_0_57525 : AO1
      port map(A => \Sensors_0_acc_z[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74829, Y => HIEFFPLA_NET_0_75020);
    
    \I2C_PassThrough_0/cnt[1]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73504, CLK => CLKINT_0_Y_0, Q
         => \I2C_PassThrough_0/cnt[1]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/we\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_72433, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72432, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_we\);
    
    HIEFFPLA_INST_0_64545 : NAND2B
      port map(A => \General_Controller_0/uc_tx_state[6]_net_1\, 
        B => \General_Controller_0/uc_tx_state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73603);
    
    HIEFFPLA_INST_0_71127 : AOI1
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        B => \Sensors_0_acc_y[4]\, C => HIEFFPLA_NET_0_71978, Y
         => HIEFFPLA_NET_0_74971);
    
    HIEFFPLA_INST_0_66248 : MX2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G3[1]_net_1\, B
         => \Science_0/ADC_READ_0_G3[1]\, S => 
        \Science_0/SET_LP_GAIN_0/state[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73168);
    
    HIEFFPLA_INST_0_63265 : AO1
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, C => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73796);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[3]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72767, Q => 
        \Sensors_0_acc_y[3]\);
    
    HIEFFPLA_INST_0_66156 : MX2B
      port map(A => \Science_0/DAC_SET_0/vector[1]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73194);
    
    HIEFFPLA_INST_0_58696 : AOI1
      port map(A => HIEFFPLA_NET_0_74517, B => 
        HIEFFPLA_NET_0_74645, C => HIEFFPLA_NET_0_74684, Y => 
        HIEFFPLA_NET_0_74702);
    
    \GS_Readout_0/subState[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74354, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/subState[1]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRY[8]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75297, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[8]\\\\\);
    
    \General_Controller_0/state_seconds[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74227, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[1]_net_1\);
    
    HIEFFPLA_INST_0_68805 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, B
         => HIEFFPLA_NET_0_72479, C => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_72553);
    
    HIEFFPLA_INST_0_58638 : AO1D
      port map(A => HIEFFPLA_NET_0_74705, B => 
        HIEFFPLA_NET_0_74655, C => HIEFFPLA_NET_0_74687, Y => 
        HIEFFPLA_NET_0_74715);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/data_out_1[6]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_72550, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72547, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[6]\);
    
    HIEFFPLA_INST_0_57519 : AO1B
      port map(A => \Sensors_0_mag_z[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75021, Y => HIEFFPLA_NET_0_75022);
    
    HIEFFPLA_INST_0_69686 : OA1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\, 
        B => HIEFFPLA_NET_0_72427, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72329);
    
    HIEFFPLA_INST_0_56025 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[10]\\\\\, B
         => HIEFFPLA_NET_0_75295, Y => HIEFFPLA_NET_0_75366);
    
    HIEFFPLA_INST_0_66061 : OR2A
      port map(A => \Science_0/DAC_SET_0/cnt[4]_net_1\, B => 
        HIEFFPLA_NET_0_73221, Y => HIEFFPLA_NET_0_73222);
    
    HIEFFPLA_INST_0_57840 : AOI1
      port map(A => \Sensors_0_acc_time[19]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74928, Y => HIEFFPLA_NET_0_74929);
    
    HIEFFPLA_INST_0_56448 : MX2
      port map(A => \FMC_DA_c[7]\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[7]\\\\\, S => 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\, Y => 
        HIEFFPLA_NET_0_75280);
    
    HIEFFPLA_INST_0_70413 : XOR2
      port map(A => HIEFFPLA_NET_0_72158, B => 
        \Timekeeper_0_microseconds[19]\, Y => 
        HIEFFPLA_NET_0_72141);
    
    HIEFFPLA_INST_0_55747 : AO1
      port map(A => HIEFFPLA_NET_0_75431, B => 
        HIEFFPLA_NET_0_75469, C => HIEFFPLA_NET_0_75429, Y => 
        HIEFFPLA_NET_0_75433);
    
    HIEFFPLA_INST_0_55477 : AXOI7
      port map(A => \Communications_0/UART_0/tx_state[0]_net_1\, 
        B => \Communications_0/UART_0/tx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_75528, Y => HIEFFPLA_NET_0_75502);
    
    HIEFFPLA_INST_0_70598 : AND3
      port map(A => \Timing_0/m_time[0]_net_1\, B => 
        HIEFFPLA_NET_0_72083, C => \Timing_0/m_time[1]_net_1\, Y
         => HIEFFPLA_NET_0_72069);
    
    HIEFFPLA_INST_0_67433 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, 
        Y => HIEFFPLA_NET_0_72882);
    
    HIEFFPLA_INST_0_61036 : AO1A
      port map(A => HIEFFPLA_NET_0_74249, B => 
        \General_Controller_0/flight_state[2]_net_1\, C => 
        HIEFFPLA_NET_0_74285, Y => HIEFFPLA_NET_0_74290);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/temp[7]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72555, Q => 
        \Sensors_0_gyro_temp[7]\);
    
    HIEFFPLA_INST_0_65151 : NAND2
      port map(A => \Sensors_0_pressure_raw[6]\, B => 
        \Sensors_0_pressure_raw[4]\, Y => HIEFFPLA_NET_0_73457);
    
    HIEFFPLA_INST_0_59550 : AO1
      port map(A => HIEFFPLA_NET_0_74429, B => 
        HIEFFPLA_NET_0_74341, C => HIEFFPLA_NET_0_74505, Y => 
        HIEFFPLA_NET_0_74539);
    
    HIEFFPLA_INST_0_66516 : NOR3B
      port map(A => HIEFFPLA_NET_0_73103, B => 
        HIEFFPLA_NET_0_73144, C => HIEFFPLA_NET_0_73146, Y => 
        HIEFFPLA_NET_0_73104);
    
    \General_Controller_0/constant_bias_probe_id[0]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73923, Q => 
        \General_Controller_0/constant_bias_probe_id[0]_net_1\);
    
    HIEFFPLA_INST_0_57644 : AOI1
      port map(A => \Science_0_exp_packet_0[33]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74982, Y => HIEFFPLA_NET_0_74983);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[4]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[4]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[4]\);
    
    \Science_0/ADC_READ_0/data_b[5]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[4]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[5]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_0[12]\ : DFN0E0P1
      port map(D => HIEFFPLA_NET_0_75241, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\);
    
    HIEFFPLA_INST_0_56960 : MX2
      port map(A => HIEFFPLA_NET_0_74970, B => 
        HIEFFPLA_NET_0_74900, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75190);
    
    HIEFFPLA_INST_0_69173 : NOR3B
      port map(A => HIEFFPLA_NET_0_72539, B => 
        HIEFFPLA_NET_0_72455, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, Y
         => HIEFFPLA_NET_0_72456);
    
    HIEFFPLA_INST_0_68451 : AO1
      port map(A => HIEFFPLA_NET_0_72645, B => 
        HIEFFPLA_NET_0_72626, C => HIEFFPLA_NET_0_72658, Y => 
        HIEFFPLA_NET_0_72647);
    
    HIEFFPLA_INST_0_61991 : AOI1C
      port map(A => HIEFFPLA_NET_0_74081, B => 
        HIEFFPLA_NET_0_74104, C => HIEFFPLA_NET_0_73889, Y => 
        HIEFFPLA_NET_0_74079);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72862, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\);
    
    HIEFFPLA_INST_0_67468 : NOR3B
      port map(A => HIEFFPLA_NET_0_72919, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, C
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72871);
    
    HIEFFPLA_INST_0_64825 : AX1C
      port map(A => HIEFFPLA_NET_0_73532, B => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, C => 
        \General_Controller_0/uc_tx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73530);
    
    \Science_0/ADC_READ_0/state[0]\ : DFN1C1
      port map(D => \Science_0/ADC_READ_0/state[1]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => 
        \Science_0/ADC_READ_0/state[0]_net_1\);
    
    HIEFFPLA_INST_0_56555 : OA1C
      port map(A => HIEFFPLA_NET_0_75241, B => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, C => 
        HIEFFPLA_NET_0_75239, Y => HIEFFPLA_NET_0_75240);
    
    HIEFFPLA_INST_0_69855 : AOI1C
      port map(A => \Sensors_0/Pressure_Sensor_0/state[8]\, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_num_bytes[1]\, 
        C => HIEFFPLA_NET_0_72288, Y => HIEFFPLA_NET_0_72290);
    
    HIEFFPLA_INST_0_62848 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[1]_net_1\, 
        B => \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        \General_Controller_0/uc_rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73883);
    
    HIEFFPLA_INST_0_62548 : AX1A
      port map(A => HIEFFPLA_NET_0_74084, B => 
        \General_Controller_0/uc_rx_byte[1]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73959);
    
    HIEFFPLA_INST_0_58314 : AO1
      port map(A => \Sensors_0_acc_y[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74803, Y => HIEFFPLA_NET_0_74804);
    
    HIEFFPLA_INST_0_68967 : AND3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, B
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_72514, Y => HIEFFPLA_NET_0_72511);
    
    HIEFFPLA_INST_0_66978 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[1]\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        C => HIEFFPLA_NET_0_72978, Y => HIEFFPLA_NET_0_72992);
    
    HIEFFPLA_INST_0_62862 : NOR3B
      port map(A => HIEFFPLA_NET_0_73921, B => 
        \General_Controller_0/uc_rx_state[0]_net_1\, C => 
        HIEFFPLA_NET_0_73811, Y => HIEFFPLA_NET_0_73879);
    
    \ClockDivs_0/cnt_800kHz[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75633, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \ClockDivs_0/cnt_800kHz[4]_net_1\);
    
    HIEFFPLA_INST_0_66118 : NOR2A
      port map(A => \Science_0/DAC_SET_0/vector[9]_net_1\, B => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73203);
    
    HIEFFPLA_INST_0_63199 : NOR2A
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73809);
    
    HIEFFPLA_INST_0_68798 : OR2A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, B
         => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, Y => 
        HIEFFPLA_NET_0_72556);
    
    \General_Controller_0/gs_id[6]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73922, Q => 
        \General_Controller_0_gs_id[6]\);
    
    HIEFFPLA_INST_0_70738 : AND3
      port map(A => \Timing_0/s_count[0]_net_1\, B => 
        HIEFFPLA_NET_0_72082, C => HIEFFPLA_NET_0_72081, Y => 
        HIEFFPLA_NET_0_72026);
    
    \Science_0/ADC_READ_0/data_a[2]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[1]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[2]_net_1\);
    
    \LDSDI_pad/U0/U0\ : IOPAD_TRI
      port map(D => \LDSDI_pad/U0/NET1\, E => \LDSDI_pad/U0/NET2\, 
        PAD => LDSDI);
    
    HIEFFPLA_INST_0_67592 : AO1E
      port map(A => HIEFFPLA_NET_0_72947, B => 
        HIEFFPLA_NET_0_72946, C => HIEFFPLA_NET_0_72957, Y => 
        HIEFFPLA_NET_0_72846);
    
    HIEFFPLA_INST_0_69590 : OR2A
      port map(A => HIEFFPLA_NET_0_72384, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_net_1\, 
        Y => HIEFFPLA_NET_0_72356);
    
    HIEFFPLA_INST_0_67547 : NAND3A
      port map(A => HIEFFPLA_NET_0_72792, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, C
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72855);
    
    HIEFFPLA_INST_0_61078 : NAND3
      port map(A => \Timekeeper_0_milliseconds[7]\, B => 
        \Timekeeper_0_milliseconds[9]\, C => 
        \Timekeeper_0_milliseconds[8]\, Y => HIEFFPLA_NET_0_74283);
    
    HIEFFPLA_INST_0_58656 : NOR2A
      port map(A => HIEFFPLA_NET_0_74484, B => 
        \General_Controller_0_gs_id[5]\, Y => 
        HIEFFPLA_NET_0_74711);
    
    \General_Controller_0/sweep_table_sample_skip[5]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[5]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[5]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[9]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72484, Q => 
        \Sensors_0_gyro_y[9]\);
    
    HIEFFPLA_INST_0_58587 : AX1C
      port map(A => HIEFFPLA_NET_0_74733, B => 
        \Eject_Signal_Debounce_0/ms_cnt[1]_net_1\, C => 
        \Eject_Signal_Debounce_0/ms_cnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74728);
    
    HIEFFPLA_INST_0_59347 : MX2
      port map(A => HIEFFPLA_NET_0_74526, B => 
        HIEFFPLA_NET_0_74578, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74565);
    
    HIEFFPLA_INST_0_65752 : AX1C
      port map(A => \Science_0/ADC_READ_0/cnt[0]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73289);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/we\ : 
        DFN1E0C1
      port map(D => \Sensors_0/Accelerometer_0/state_0[8]\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72710, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_we\);
    
    HIEFFPLA_INST_0_62126 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => HIEFFPLA_NET_0_73916, C => HIEFFPLA_NET_0_73890, Y
         => HIEFFPLA_NET_0_74046);
    
    HIEFFPLA_INST_0_58760 : NAND3C
      port map(A => HIEFFPLA_NET_0_74681, B => 
        HIEFFPLA_NET_0_74678, C => HIEFFPLA_NET_0_74676, Y => 
        HIEFFPLA_NET_0_74691);
    
    HIEFFPLA_INST_0_66686 : AND2B
      port map(A => ACCE_SCL_c, B => 
        \Sensors_0/Accelerometer_0/state_0[8]\, Y => 
        HIEFFPLA_NET_0_73065);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[8]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[8]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[8]\);
    
    HIEFFPLA_INST_0_68797 : NAND2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, B
         => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, Y => 
        HIEFFPLA_NET_0_72557);
    
    HIEFFPLA_INST_0_66283 : NAND2
      port map(A => HIEFFPLA_NET_0_73171, B => 
        \Science_0/SET_LP_GAIN_0/state[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73156);
    
    HIEFFPLA_INST_0_55376 : XA1C
      port map(A => HIEFFPLA_NET_0_75501, B => 
        \Communications_0/UART_0/tx_clk_count[0]_net_1\, C => 
        HIEFFPLA_NET_0_75527, Y => HIEFFPLA_NET_0_75526);
    
    HIEFFPLA_INST_0_58363 : AND2
      port map(A => \Sensors_0_mag_y[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        Y => HIEFFPLA_NET_0_74791);
    
    \Science_0/ADC_READ_0/exp_packet_1[33]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[17]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[33]\);
    
    HIEFFPLA_INST_0_68367 : AND2
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[0]_net_1\, B
         => \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72669);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[9]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72553, Q => 
        \Sensors_0_gyro_x[9]\);
    
    HIEFFPLA_INST_0_59367 : MX2
      port map(A => HIEFFPLA_NET_0_74492, B => 
        HIEFFPLA_NET_0_74375, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74563);
    
    HIEFFPLA_INST_0_68196 : NOR3B
      port map(A => HIEFFPLA_NET_0_72708, B => 
        HIEFFPLA_NET_0_72912, C => HIEFFPLA_NET_0_72893, Y => 
        HIEFFPLA_NET_0_72709);
    
    \Communications_0/UART_1/recv[1]\ : DFN1E1C1
      port map(D => \Communications_0/UART_1/rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75441, Q => \Communications_0_uc_recv[1]\);
    
    HIEFFPLA_INST_0_64509 : AND3B
      port map(A => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, B => 
        HIEFFPLA_NET_0_73552, C => 
        \General_Controller_0/uc_tx_state[12]_net_1\, Y => 
        HIEFFPLA_NET_0_73610);
    
    HIEFFPLA_INST_0_67138 : AND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[6]_net_1\, 
        Y => HIEFFPLA_NET_0_72955);
    
    HIEFFPLA_INST_0_70581 : NOR2A
      port map(A => HIEFFPLA_NET_0_72072, B => 
        HIEFFPLA_NET_0_72083, Y => HIEFFPLA_NET_0_72073);
    
    HIEFFPLA_INST_0_66066 : AND2B
      port map(A => \Science_0/DAC_SET_0/cnt[2]_net_1\, B => 
        \Science_0/DAC_SET_0/cnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73220);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[13]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[13]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[13]\);
    
    HIEFFPLA_INST_0_64494 : NOR2A
      port map(A => \General_Controller_0/uc_tx_state[14]_net_1\, 
        B => \General_Controller_0/uc_tx_substate[1]_net_1\, Y
         => HIEFFPLA_NET_0_73615);
    
    HIEFFPLA_INST_0_65675 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt4dn[6]_net_1\, B => 
        HIEFFPLA_NET_0_73327, C => HIEFFPLA_NET_0_73274, Y => 
        HIEFFPLA_NET_0_73312);
    
    HIEFFPLA_INST_0_59087 : OA1A
      port map(A => HIEFFPLA_NET_0_74432, B => 
        HIEFFPLA_NET_0_74725, C => \GS_Readout_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_74617);
    
    HIEFFPLA_INST_0_58619 : AND3
      port map(A => HIEFFPLA_NET_0_74724, B => 
        HIEFFPLA_NET_0_74723, C => HIEFFPLA_NET_0_74721, Y => 
        HIEFFPLA_NET_0_74718);
    
    \General_Controller_0/sweep_table_points[15]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[15]_net_1\);
    
    \Eject_Signal_Debounce_0/ms_cnt[0]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74747, CLK => CLKINT_0_Y_0, Q
         => \Eject_Signal_Debounce_0/ms_cnt[0]_net_1\);
    
    \Communications_0/UART_0/tx_clk_count[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75526, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_clk_count[0]_net_1\);
    
    HIEFFPLA_INST_0_58003 : AO1
      port map(A => \Science_0_exp_packet_0[55]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75122, Y => HIEFFPLA_NET_0_74882);
    
    HIEFFPLA_INST_0_68349 : AND3A
      port map(A => HIEFFPLA_NET_0_72674, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, C => 
        GYRO_SCL_c, Y => HIEFFPLA_NET_0_72675);
    
    \Timing_0/s_time[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72047, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \s_clks_net_0[18]\);
    
    \Science_0/SWEEP_SPIDER2_0/update\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73151, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Science_0/SWEEP_SPIDER2_0_SET\);
    
    HIEFFPLA_INST_0_60977 : AOI1D
      port map(A => \Timekeeper_0_milliseconds[3]\, B => 
        \Timekeeper_0_milliseconds[4]\, C => 
        \General_Controller_0/flight_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74305);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_2\ : 
        DFN0E0P1
      port map(D => HIEFFPLA_NET_0_72359, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72384, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_2_net_1\);
    
    \Pressure_Signal_Debounce_0/ms_cnt[6]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73488, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[6]_net_1\);
    
    \General_Controller_0/constant_bias_voltage_0[9]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[9]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72219, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]_net_1\);
    
    HIEFFPLA_INST_0_61186 : NAND3C
      port map(A => 
        \General_Controller_0/state_seconds[12]_net_1\, B => 
        \General_Controller_0/state_seconds[14]_net_1\, C => 
        \General_Controller_0/state_seconds[17]_net_1\, Y => 
        HIEFFPLA_NET_0_74256);
    
    HIEFFPLA_INST_0_62043 : NAND3C
      port map(A => HIEFFPLA_NET_0_73953, B => 
        HIEFFPLA_NET_0_73898, C => HIEFFPLA_NET_0_74067, Y => 
        HIEFFPLA_NET_0_74064);
    
    HIEFFPLA_INST_0_55854 : AXOI7
      port map(A => HIEFFPLA_NET_0_75420, B => 
        HIEFFPLA_NET_0_75386, C => 
        \Communications_0/UART_1/tx_clk_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75411);
    
    HIEFFPLA_INST_0_71130 : AOI1D
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => \Sensors_0_acc_temp[4]\, Y => HIEFFPLA_NET_0_71977);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72769, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\);
    
    HIEFFPLA_INST_0_70427 : AX1C
      port map(A => \Timekeeper_0_microseconds[0]\, B => 
        \Timekeeper_0_microseconds[1]\, C => 
        \Timekeeper_0_microseconds[2]\, Y => HIEFFPLA_NET_0_72135);
    
    HIEFFPLA_INST_0_69303 : NAND3C
      port map(A => HIEFFPLA_NET_0_72426, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\, 
        C => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72424);
    
    HIEFFPLA_INST_0_66399 : AX1B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        C => HIEFFPLA_NET_0_73126, Y => HIEFFPLA_NET_0_73129);
    
    HIEFFPLA_INST_0_58693 : NAND3B
      port map(A => HIEFFPLA_NET_0_74672, B => 
        HIEFFPLA_NET_0_74679, C => HIEFFPLA_NET_0_74702, Y => 
        HIEFFPLA_NET_0_74703);
    
    HIEFFPLA_INST_0_67925 : NOR3A
      port map(A => HIEFFPLA_NET_0_72780, B => 
        HIEFFPLA_NET_0_72880, C => HIEFFPLA_NET_0_72896, Y => 
        HIEFFPLA_NET_0_72772);
    
    \General_Controller_0/st_wdata[15]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[15]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[15]\);
    
    HIEFFPLA_INST_0_58660 : AO1
      port map(A => \General_Controller_0_gs_id[6]\, B => 
        HIEFFPLA_NET_0_74484, C => HIEFFPLA_NET_0_74709, Y => 
        HIEFFPLA_NET_0_74710);
    
    HIEFFPLA_INST_0_56466 : XNOR2
      port map(A => HIEFFPLA_NET_0_75321, B => 
        HIEFFPLA_NET_0_75318, Y => HIEFFPLA_NET_0_75273);
    
    HIEFFPLA_INST_0_70082 : OR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72226);
    
    HIEFFPLA_INST_0_58970 : OA1A
      port map(A => HIEFFPLA_NET_0_74521, B => 
        HIEFFPLA_NET_0_74457, C => \GS_Readout_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_74646);
    
    HIEFFPLA_INST_0_66864 : AND3A
      port map(A => HIEFFPLA_NET_0_73017, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73018);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1E1C0_data_out[4]\\\\/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75283, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \FMC_DA_c[4]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/data_out_1[3]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_72554, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72547, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[3]\);
    
    HIEFFPLA_INST_0_61096 : NOR3A
      port map(A => HIEFFPLA_NET_0_74277, B => 
        \Timekeeper_0_milliseconds[16]\, C => 
        \Timekeeper_0_milliseconds[15]\, Y => 
        HIEFFPLA_NET_0_74278);
    
    HIEFFPLA_INST_0_55588 : OR3B
      port map(A => HIEFFPLA_NET_0_75472, B => 
        \Communications_0/UART_1/rx_clk_count_c0\, C => 
        \Communications_0/UART_1/rx_clk_count[25]_net_1\, Y => 
        HIEFFPLA_NET_0_75473);
    
    HIEFFPLA_INST_0_60894 : OR3A
      port map(A => \General_Controller_0/command[4]_net_1\, B
         => \General_Controller_0/command[2]_net_1\, C => 
        \General_Controller_0/command[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74327);
    
    HIEFFPLA_INST_0_58595 : NAND3
      port map(A => \Eject_Signal_Debounce_0/ms_cnt[3]_net_1\, B
         => HIEFFPLA_NET_0_74733, C => 
        \Eject_Signal_Debounce_0/ms_cnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74726);
    
    HIEFFPLA_INST_0_67205 : OA1A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        C => HIEFFPLA_NET_0_72929, Y => HIEFFPLA_NET_0_72940);
    
    HIEFFPLA_INST_0_55192 : NAND2
      port map(A => \Communications_0/UART_0/rx_count[1]_net_1\, 
        B => \Communications_0/UART_0/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75562);
    
    HIEFFPLA_INST_0_69008 : AND3
      port map(A => HIEFFPLA_NET_0_72540, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        C => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72499);
    
    HIEFFPLA_INST_0_62154 : AOI1D
      port map(A => HIEFFPLA_NET_0_73783, B => 
        HIEFFPLA_NET_0_73930, C => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74041);
    
    HIEFFPLA_INST_0_61220 : OR2A
      port map(A => 
        \General_Controller_0/state_seconds[12]_net_1\, B => 
        HIEFFPLA_NET_0_74251, Y => HIEFFPLA_NET_0_74246);
    
    HIEFFPLA_INST_0_56303 : XOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, B
         => HIEFFPLA_NET_0_75349, C => HIEFFPLA_NET_0_75260, Y
         => HIEFFPLA_NET_0_75313);
    
    HIEFFPLA_INST_0_55102 : NAND3
      port map(A => HIEFFPLA_NET_0_75595, B => 
        \Communications_0/UART_0/rx_clk_count_c0\, C => 
        \Communications_0/UART_0/rx_clk_count[28]_net_1\, Y => 
        HIEFFPLA_NET_0_75590);
    
    HIEFFPLA_INST_0_61468 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[51]\, B => 
        \Timekeeper_0_milliseconds[11]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74195);
    
    HIEFFPLA_INST_0_59053 : AND3C
      port map(A => HIEFFPLA_NET_0_74644, B => 
        HIEFFPLA_NET_0_74642, C => HIEFFPLA_NET_0_74656, Y => 
        HIEFFPLA_NET_0_74625);
    
    \Data_Saving_0/Packet_Saver_0/acc_flag\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_75240, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => 
        General_Controller_0_en_data_saving, Q => 
        \Data_Saving_0/Packet_Saver_0/acc_flag_net_1\);
    
    \FMC_DA_pad[6]/U0/U0\ : IOPAD_TRI
      port map(D => \FMC_DA_pad[6]/U0/NET1\, E => 
        \FMC_DA_pad[6]/U0/NET2\, PAD => FMC_DA(6));
    
    HIEFFPLA_INST_0_68565 : AND2B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, B => 
        \Sensors_0/Gyro_0/state[8]\, Y => HIEFFPLA_NET_0_72616);
    
    HIEFFPLA_INST_0_88375 : XA1A
      port map(A => HIEFFPLA_NET_0_88382, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[9]\\\\\, C => 
        HIEFFPLA_NET_0_75291, Y => HIEFFPLA_NET_0_89694);
    
    \General_Controller_0/sweep_table_read_value[13]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74166, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[13]_net_1\);
    
    HIEFFPLA_INST_0_55212 : OA1A
      port map(A => HIEFFPLA_NET_0_75562, B => 
        \Communications_0/UART_0/rx_count[2]_net_1\, C => 
        \Communications_0/UART_0/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75559);
    
    \Science_0/ADC_READ_0/cnt4dn[3]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73315, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4dn[3]_net_1\);
    
    HIEFFPLA_INST_0_61663 : MX2
      port map(A => \SweepTable_0_RD[15]\, B => 
        \SweepTable_1_RD[15]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74164);
    
    HIEFFPLA_INST_0_62480 : AND3
      port map(A => \General_Controller_0/uc_rx_state[4]_net_1\, 
        B => \General_Controller_0/uc_rx_state[3]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73974);
    
    HIEFFPLA_INST_0_68156 : NAND3C
      port map(A => HIEFFPLA_NET_0_72922, B => 
        HIEFFPLA_NET_0_72906, C => HIEFFPLA_NET_0_72719, Y => 
        HIEFFPLA_NET_0_72720);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[3]\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72405, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72352, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[3]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[1]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72482, Q => 
        \Sensors_0_gyro_y[1]\);
    
    HIEFFPLA_INST_0_71010 : AND2B
      port map(A => HIEFFPLA_NET_0_71990, B => UC_I2C4_SDA_in, Y
         => HIEFFPLA_NET_0_73510);
    
    HIEFFPLA_INST_0_57788 : AOI1
      port map(A => \Science_0_exp_packet_0[52]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74781, Y => HIEFFPLA_NET_0_74942);
    
    \Communications_0/UART_0/tx_count[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75509, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75503, Q => 
        \Communications_0/UART_0/tx_count[0]_net_1\);
    
    HIEFFPLA_INST_0_67147 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[2]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72952);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_72421, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\);
    
    HIEFFPLA_INST_0_56382 : AX1
      port map(A => HIEFFPLA_NET_0_75372, B => 
        HIEFFPLA_NET_0_75376, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[8]\\\\\, Y
         => HIEFFPLA_NET_0_75295);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[11]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72283, Q => 
        \Sensors_0_pressure_temp_raw[11]\);
    
    HIEFFPLA_INST_0_71007 : AOI1A
      port map(A => HIEFFPLA_NET_0_73439, B => 
        HIEFFPLA_NET_0_73481, C => 
        \Pressure_Signal_Debounce_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_71992);
    
    HIEFFPLA_INST_0_58943 : NAND2B
      port map(A => \GS_Readout_0/state[6]_net_1\, B => 
        \GS_Readout_0/state[7]_net_1\, Y => HIEFFPLA_NET_0_74653);
    
    \General_Controller_0/st_wdata[9]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[9]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[9]\);
    
    HIEFFPLA_INST_0_67986 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => HIEFFPLA_NET_0_72737, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72761);
    
    HIEFFPLA_INST_0_58785 : AND2
      port map(A => HIEFFPLA_NET_0_74397, B => 
        HIEFFPLA_NET_0_74645, Y => HIEFFPLA_NET_0_74685);
    
    HIEFFPLA_INST_0_65326 : AND2
      port map(A => \Science_0/ADC_READ_0/cnt1dn[0]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt1dn[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73409);
    
    \General_Controller_0/constant_bias_voltage_1[9]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[9]_net_1\);
    
    \General_Controller_0/status_bits_1[45]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74201, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[45]\);
    
    \Communications_0/UART_0/tx_state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75500, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_state[0]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRY[9]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75306, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[9]\\\\\);
    
    HIEFFPLA_INST_0_65903 : AND2B
      port map(A => \Science_0/ADC_READ_0_G1[0]\, B => 
        \Science_0/ADC_READ_0_G1[1]\, Y => HIEFFPLA_NET_0_73261);
    
    HIEFFPLA_INST_0_68723 : AO1A
      port map(A => HIEFFPLA_NET_0_72689, B => 
        HIEFFPLA_NET_0_72631, C => HIEFFPLA_NET_0_72576, Y => 
        HIEFFPLA_NET_0_72578);
    
    HIEFFPLA_INST_0_66007 : OA1A
      port map(A => HIEFFPLA_NET_0_73299, B => 
        HIEFFPLA_NET_0_73296, C => 
        \Science_0/ADC_READ_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73239);
    
    \General_Controller_0/sweep_table_step_id[4]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73926, Q => 
        \General_Controller_0/sweep_table_step_id[4]_net_1\);
    
    HIEFFPLA_INST_0_62770 : AND3
      port map(A => HIEFFPLA_NET_0_73883, B => 
        HIEFFPLA_NET_0_73780, C => HIEFFPLA_NET_0_73888, Y => 
        HIEFFPLA_NET_0_73910);
    
    HIEFFPLA_INST_0_59605 : MX2
      port map(A => HIEFFPLA_NET_0_74453, B => 
        HIEFFPLA_NET_0_74381, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74532);
    
    \Science_0/ADC_READ_0/cnt2up[4]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73360, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2up[4]_net_1\);
    
    HIEFFPLA_INST_0_61894 : NOR3B
      port map(A => \General_Controller_0/uc_rx_byte[2]_net_1\, B
         => \General_Controller_0/uc_rx_substate[2]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74106);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[8]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72490, Q => 
        \ch3_data_net_0[4]\);
    
    HIEFFPLA_INST_0_66078 : XNOR2
      port map(A => HIEFFPLA_NET_0_73225, B => 
        \Science_0/DAC_SET_0/cnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73216);
    
    HIEFFPLA_INST_0_60851 : XNOR2
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74342);
    
    HIEFFPLA_INST_0_62468 : NAND3C
      port map(A => HIEFFPLA_NET_0_73868, B => 
        HIEFFPLA_NET_0_74008, C => HIEFFPLA_NET_0_74097, Y => 
        HIEFFPLA_NET_0_73976);
    
    HIEFFPLA_INST_0_58809 : AO1
      port map(A => HIEFFPLA_NET_0_74421, B => 
        HIEFFPLA_NET_0_74633, C => HIEFFPLA_NET_0_74664, Y => 
        HIEFFPLA_NET_0_74681);
    
    HIEFFPLA_INST_0_58919 : AO1C
      port map(A => HIEFFPLA_NET_0_74671, B => 
        HIEFFPLA_NET_0_74661, C => HIEFFPLA_NET_0_74658, Y => 
        HIEFFPLA_NET_0_74659);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[0]\ : 
        DFN0C1
      port map(D => HIEFFPLA_NET_0_72408, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[0]_net_1\);
    
    HIEFFPLA_INST_0_63396 : MX2
      port map(A => HIEFFPLA_NET_0_73759, B => 
        HIEFFPLA_NET_0_73694, S => HIEFFPLA_NET_0_73608, Y => 
        HIEFFPLA_NET_0_73767);
    
    \Sensors_0/Gyro_0/I2C_Master_0/data_out[0]\ : DFN0E1C1
      port map(D => GYRO_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72683, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[0]\);
    
    HIEFFPLA_INST_0_67848 : AND3
      port map(A => HIEFFPLA_NET_0_72809, B => 
        HIEFFPLA_NET_0_72872, C => HIEFFPLA_NET_0_72911, Y => 
        HIEFFPLA_NET_0_72788);
    
    HIEFFPLA_INST_0_66000 : OR2A
      port map(A => \Science_0/ADC_READ_0/newflag_net_1\, B => 
        CLKINT_1_Y, Y => HIEFFPLA_NET_0_73243);
    
    HIEFFPLA_INST_0_64695 : NOR2A
      port map(A => Communications_0_uc_tx_rdy, B => 
        HIEFFPLA_NET_0_73558, Y => HIEFFPLA_NET_0_73561);
    
    HIEFFPLA_INST_0_70716 : AND3
      port map(A => \Timing_0/s_time[1]_net_1\, B => 
        \Timing_0/s_time[0]_net_1\, C => HIEFFPLA_NET_0_72058, Y
         => HIEFFPLA_NET_0_72033);
    
    HIEFFPLA_INST_0_57798 : AOI1
      port map(A => \Science_0_exp_packet_0[53]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74813, Y => HIEFFPLA_NET_0_74939);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/i2c_repeat_start\ : 
        DFN1E0C1
      port map(D => HIEFFPLA_NET_0_72492, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72562, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_i2c_repeat_start\);
    
    HIEFFPLA_INST_0_68076 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72737);
    
    HIEFFPLA_INST_0_62593 : NOR3B
      port map(A => HIEFFPLA_NET_0_73949, B => 
        HIEFFPLA_NET_0_73901, C => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73950);
    
    \Data_Saving_0/Packet_Saver_0/packet_select[12]\ : DFN0E0P1
      port map(D => HIEFFPLA_NET_0_75241, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\);
    
    HIEFFPLA_INST_0_67996 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72758);
    
    HIEFFPLA_INST_0_63848 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[4]_net_1\, B
         => 
        \General_Controller_0/sweep_table_sample_skip[4]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73701);
    
    HIEFFPLA_INST_0_63548 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[10]_net_1\, B
         => \General_Controller_0/sweep_table_points[10]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73751);
    
    HIEFFPLA_INST_0_57267 : AND2
      port map(A => \Sensors_0_acc_y[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        Y => HIEFFPLA_NET_0_75103);
    
    HIEFFPLA_INST_0_65147 : NAND3
      port map(A => HIEFFPLA_NET_0_73458, B => 
        \Sensors_0_pressure_raw[15]\, C => 
        \Sensors_0_pressure_raw[17]\, Y => HIEFFPLA_NET_0_73459);
    
    HIEFFPLA_INST_0_62791 : NOR3A
      port map(A => HIEFFPLA_NET_0_74063, B => 
        HIEFFPLA_NET_0_74068, C => HIEFFPLA_NET_0_73902, Y => 
        HIEFFPLA_NET_0_73903);
    
    HIEFFPLA_INST_0_55485 : AO1
      port map(A => HIEFFPLA_NET_0_75512, B => 
        \Communications_0/UART_0/tx_count[1]_net_1\, C => 
        HIEFFPLA_NET_0_75498, Y => HIEFFPLA_NET_0_75500);
    
    \Science_0/ADC_READ_0/chan4_data[4]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[4]\);
    
    HIEFFPLA_INST_0_68319 : AND3
      port map(A => HIEFFPLA_NET_0_72702, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, C => 
        GYRO_SCL_c, Y => HIEFFPLA_NET_0_72683);
    
    HIEFFPLA_INST_0_64673 : AND2
      port map(A => 
        \General_Controller_0/uc_tx_nextstate[4]_net_1\, B => 
        HIEFFPLA_NET_0_73584, Y => HIEFFPLA_NET_0_73569);
    
    HIEFFPLA_INST_0_58823 : AND2
      port map(A => HIEFFPLA_NET_0_74521, B => 
        HIEFFPLA_NET_0_74646, Y => HIEFFPLA_NET_0_74679);
    
    HIEFFPLA_INST_0_58555 : XA1A
      port map(A => \Eject_Signal_Debounce_0/state[0]_net_1\, B
         => HIEFFPLA_NET_0_74736, C => HIEFFPLA_NET_0_74749, Y
         => HIEFFPLA_NET_0_74735);
    
    HIEFFPLA_INST_0_56513 : AX1C
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, B
         => HIEFFPLA_NET_0_75349, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\, Y
         => HIEFFPLA_NET_0_75258);
    
    HIEFFPLA_INST_0_60575 : MX2
      port map(A => \Science_0_chan6_data[4]\, B => 
        \Science_0_chan6_data[8]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74393);
    
    HIEFFPLA_INST_0_55558 : NOR3B
      port map(A => HIEFFPLA_NET_0_75478, B => 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\, C => 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\, Y => 
        HIEFFPLA_NET_0_75481);
    
    \General_Controller_0/sweep_table_sweep_cnt[9]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74129, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[9]_net_1\);
    
    HIEFFPLA_INST_0_68381 : AND2B
      port map(A => HIEFFPLA_NET_0_72689, B => GYRO_SCL_c, Y => 
        HIEFFPLA_NET_0_72663);
    
    HIEFFPLA_INST_0_71368 : OA1A
      port map(A => HIEFFPLA_NET_0_72745, B => 
        HIEFFPLA_NET_0_72752, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_71969);
    
    HIEFFPLA_INST_0_65091 : MX2A
      port map(A => HIEFFPLA_NET_0_73472, B => 
        HIEFFPLA_NET_0_73481, S => 
        \Pressure_Signal_Debounce_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73473);
    
    HIEFFPLA_INST_0_67285 : AND3C
      port map(A => HIEFFPLA_NET_0_72927, B => 
        HIEFFPLA_NET_0_72759, C => HIEFFPLA_NET_0_72898, Y => 
        HIEFFPLA_NET_0_72917);
    
    HIEFFPLA_INST_0_60410 : MX2
      port map(A => HIEFFPLA_NET_0_74422, B => 
        HIEFFPLA_NET_0_74540, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74419);
    
    \Communications_0/UART_0/rx_byte[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75380, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75612, Q => 
        \Communications_0/UART_0/rx_byte[0]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[4]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72482, Q => 
        \Sensors_0_gyro_y[4]\);
    
    HIEFFPLA_INST_0_55145 : XA1B
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[24]_net_1\, B => 
        HIEFFPLA_NET_0_75598, C => HIEFFPLA_NET_0_75567, Y => 
        HIEFFPLA_NET_0_75575);
    
    HIEFFPLA_INST_0_55961 : AX1
      port map(A => HIEFFPLA_NET_0_75420, B => 
        \Communications_0/UART_1/tx_state[0]_net_1\, C => 
        \Communications_0/UART_1/tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75383);
    
    HIEFFPLA_INST_0_70138 : OA1C
      port map(A => HIEFFPLA_NET_0_72267, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]_net_1\, 
        C => HIEFFPLA_NET_0_72205, Y => HIEFFPLA_NET_0_72211);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[6]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[6]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[6]\);
    
    HIEFFPLA_INST_0_67166 : AND3
      port map(A => HIEFFPLA_NET_0_72955, B => 
        HIEFFPLA_NET_0_72960, C => HIEFFPLA_NET_0_72950, Y => 
        HIEFFPLA_NET_0_72947);
    
    HIEFFPLA_INST_0_58767 : AO1
      port map(A => HIEFFPLA_NET_0_74646, B => 
        HIEFFPLA_NET_0_74510, C => HIEFFPLA_NET_0_74689, Y => 
        HIEFFPLA_NET_0_74690);
    
    HIEFFPLA_INST_0_67503 : AND2B
      port map(A => HIEFFPLA_NET_0_72915, B => 
        HIEFFPLA_NET_0_72851, Y => HIEFFPLA_NET_0_72863);
    
    HIEFFPLA_INST_0_64759 : AO1A
      port map(A => HIEFFPLA_NET_0_73613, B => 
        HIEFFPLA_NET_0_73546, C => HIEFFPLA_NET_0_73547, Y => 
        HIEFFPLA_NET_0_73548);
    
    \General_Controller_0/command[1]\ : DFN1E1
      port map(D => \Communications_0_ext_recv[1]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74300, Q => 
        \General_Controller_0/command[1]_net_1\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_72696, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\);
    
    HIEFFPLA_INST_0_66843 : AO1D
      port map(A => HIEFFPLA_NET_0_73060, B => 
        HIEFFPLA_NET_0_73101, C => HIEFFPLA_NET_0_73018, Y => 
        HIEFFPLA_NET_0_73023);
    
    HIEFFPLA_INST_0_66151 : MX2B
      port map(A => \Science_0/DAC_SET_0/vector[0]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73195);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[8]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72753, Q => 
        \Sensors_0_acc_z[8]\);
    
    HIEFFPLA_INST_0_61779 : XOR2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[0]_net_1\, B
         => \General_Controller_0/sweep_table_sweep_cnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_74137);
    
    \Science_0/ADC_READ_0/g2i[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73260, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73420, Q => 
        \Science_0/ADC_READ_0_G2[0]\);
    
    \Timing_0/m_time[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72066, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_time[3]_net_1\);
    
    HIEFFPLA_INST_0_63836 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[2]_net_1\, B
         => 
        \General_Controller_0/sweep_table_sample_skip[2]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73703);
    
    \Sensors_0/Gyro_0/I2C_Master_0/scl_0\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_72633, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\);
    
    HIEFFPLA_INST_0_57675 : AO1B
      port map(A => \Sensors_0_acc_x[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74973, Y => HIEFFPLA_NET_0_74974);
    
    HIEFFPLA_INST_0_62452 : AND2
      port map(A => HIEFFPLA_NET_0_73972, B => 
        HIEFFPLA_NET_0_73778, Y => HIEFFPLA_NET_0_73979);
    
    HIEFFPLA_INST_0_59824 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[59]\, B => 
        \Data_Hub_Packets_0_status_packet[63]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74502);
    
    HIEFFPLA_INST_0_55529 : NOR3A
      port map(A => \Communications_0/UART_1/rx_count[0]_net_1\, 
        B => \Communications_0/UART_1/rx_count[2]_net_1\, C => 
        \Communications_0/UART_1/rx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75486);
    
    \General_Controller_0/sweep_table_write_value[14]\ : DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[14]_net_1\);
    
    HIEFFPLA_INST_0_56731 : AOI1C
      port map(A => HIEFFPLA_NET_0_75186, B => 
        HIEFFPLA_NET_0_75187, C => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75220);
    
    HIEFFPLA_INST_0_88374 : XAI1A
      port map(A => HIEFFPLA_NET_0_75304, B => 
        HIEFFPLA_NET_0_75320, C => HIEFFPLA_NET_0_75326, Y => 
        HIEFFPLA_NET_0_88383);
    
    HIEFFPLA_INST_0_71034 : NAND3B
      port map(A => \General_Controller_0/uc_tx_state[3]_net_1\, 
        B => \General_Controller_0/uc_tx_state[0]_net_1\, C => 
        HIEFFPLA_NET_0_73596, Y => HIEFFPLA_NET_0_71986);
    
    HIEFFPLA_INST_0_62233 : XA1
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[1]_net_1\, C => 
        HIEFFPLA_NET_0_73974, Y => HIEFFPLA_NET_0_74024);
    
    HIEFFPLA_INST_0_65316 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt1dn[3]_net_1\, B => 
        HIEFFPLA_NET_0_73410, C => 
        \Science_0/ADC_READ_0/cnt1dn[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73413);
    
    HIEFFPLA_INST_0_59111 : AND3
      port map(A => HIEFFPLA_NET_0_74593, B => 
        HIEFFPLA_NET_0_74723, C => HIEFFPLA_NET_0_74720, Y => 
        HIEFFPLA_NET_0_74610);
    
    HIEFFPLA_INST_0_70970 : XA1A
      port map(A => HIEFFPLA_NET_0_71998, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[3]_net_1\, 
        C => HIEFFPLA_NET_0_73063, Y => HIEFFPLA_NET_0_73136);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[1]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72919, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[1]_net_1\);
    
    HIEFFPLA_INST_0_68238 : NOR3B
      port map(A => HIEFFPLA_NET_0_72702, B => 
        HIEFFPLA_NET_0_72624, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_72698);
    
    \General_Controller_0/sweep_table_sample_skip[3]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[3]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[3]_net_1\);
    
    \GS_Readout_0/state[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74604, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/state[4]_net_1\);
    
    HIEFFPLA_INST_0_55734 : AND2B
      port map(A => HIEFFPLA_NET_0_75433, B => 
        HIEFFPLA_NET_0_75441, Y => HIEFFPLA_NET_0_75435);
    
    HIEFFPLA_INST_0_65820 : AO1A
      port map(A => HIEFFPLA_NET_0_73328, B => 
        HIEFFPLA_NET_0_73277, C => HIEFFPLA_NET_0_73422, Y => 
        HIEFFPLA_NET_0_73274);
    
    HIEFFPLA_INST_0_61345 : AX1B
      port map(A => HIEFFPLA_NET_0_74248, B => 
        HIEFFPLA_NET_0_74245, C => 
        \General_Controller_0/state_seconds[7]_net_1\, Y => 
        HIEFFPLA_NET_0_74211);
    
    HIEFFPLA_INST_0_60555 : MX2
      port map(A => \Science_0_chan3_data[10]\, B => 
        \Science_0_chan2_data[2]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74396);
    
    HIEFFPLA_INST_0_65184 : AX1C
      port map(A => HIEFFPLA_NET_0_73444, B => 
        \Pressure_Signal_Debounce_0/ms_cnt[4]_net_1\, C => 
        \Pressure_Signal_Debounce_0/ms_cnt[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73450);
    
    HIEFFPLA_INST_0_57240 : AND2B
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        Y => HIEFFPLA_NET_0_75117);
    
    HIEFFPLA_INST_0_69441 : AND3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[2]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72389);
    
    HIEFFPLA_INST_0_59238 : AOI1C
      port map(A => HIEFFPLA_NET_0_74382, B => 
        \GS_Readout_0/state[3]_net_1\, C => 
        Communications_0_ext_tx_rdy, Y => HIEFFPLA_NET_0_74581);
    
    \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]\ : DFN0E0
      port map(D => HIEFFPLA_NET_0_72666, CLK => 
        ClockDivs_0_clk_800kHz, E => HIEFFPLA_NET_0_72617, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\);
    
    \Science_0/ADC_READ_0/cnt3dn[7]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73340, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3dn[7]_net_1\);
    
    HIEFFPLA_INST_0_66752 : NAND3
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_repeat_start\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73046);
    
    HIEFFPLA_INST_0_57565 : AO1B
      port map(A => \Sensors_0_gyro_x[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75006, Y => HIEFFPLA_NET_0_75007);
    
    HIEFFPLA_INST_0_62019 : XA1B
      port map(A => 
        \General_Controller_0/uc_rx_prev_state[2]_net_1\, B => 
        \General_Controller_0/uc_rx_prev_state[3]_net_1\, C => 
        Communications_0_uc_rx_rdy, Y => HIEFFPLA_NET_0_74070);
    
    HIEFFPLA_INST_0_68189 : NOR3B
      port map(A => HIEFFPLA_NET_0_72716, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => HIEFFPLA_NET_0_72764, Y => HIEFFPLA_NET_0_72711);
    
    HIEFFPLA_INST_0_58664 : AND3C
      port map(A => HIEFFPLA_NET_0_74655, B => 
        \GS_Readout_0/state[0]_net_1\, C => HIEFFPLA_NET_0_74650, 
        Y => HIEFFPLA_NET_0_74709);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_WADDR[3]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75299, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\);
    
    HIEFFPLA_INST_0_55580 : NAND2
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[30]_net_1\, B => 
        \Communications_0/UART_1/rx_clk_count_c0\, Y => 
        HIEFFPLA_NET_0_75475);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[16]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[16]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[16]\);
    
    \General_Controller_0/sweep_table_write_value[7]\ : DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[7]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[7]_net_1\);
    
    \General_Controller_0/status_bits_1[46]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74200, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[46]\);
    
    HIEFFPLA_INST_0_63890 : MX2
      port map(A => HIEFFPLA_NET_0_73669, B => 
        HIEFFPLA_NET_0_73663, S => HIEFFPLA_NET_0_73594, Y => 
        HIEFFPLA_NET_0_73694);
    
    HIEFFPLA_INST_0_68995 : NOR3A
      port map(A => HIEFFPLA_NET_0_72508, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72504);
    
    HIEFFPLA_INST_0_66231 : MX2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G2[1]_net_1\, B
         => \Science_0/ADC_READ_0_G2[1]\, S => 
        \Science_0/SET_LP_GAIN_0/state[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73172);
    
    \Science_0/ADC_READ_0/data_b[3]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[2]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[3]_net_1\);
    
    \Science_0/ADC_READ_0/chan1_data[6]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[6]\);
    
    HIEFFPLA_INST_0_59077 : OA1A
      port map(A => HIEFFPLA_NET_0_74474, B => 
        HIEFFPLA_NET_0_74468, C => \GS_Readout_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_74620);
    
    HIEFFPLA_INST_0_58723 : NOR3B
      port map(A => HIEFFPLA_NET_0_74652, B => 
        HIEFFPLA_NET_0_74569, C => HIEFFPLA_NET_0_74574, Y => 
        HIEFFPLA_NET_0_74697);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[14]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72490, Q => 
        \ch3_data_net_0[10]\);
    
    HIEFFPLA_INST_0_55334 : MX2C
      port map(A => \Communications_0/UART_0/tx_byte[1]_net_1\, B
         => \Communications_0/UART_0/tx_byte[5]_net_1\, S => 
        \Communications_0/UART_0/tx_count[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75538);
    
    HIEFFPLA_INST_0_61768 : AX1C
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[11]_net_1\, B
         => HIEFFPLA_NET_0_74149, C => 
        \General_Controller_0/sweep_table_sweep_cnt[12]_net_1\, Y
         => HIEFFPLA_NET_0_74141);
    
    HIEFFPLA_INST_0_70432 : XOR2
      port map(A => HIEFFPLA_NET_0_72156, B => 
        \Timekeeper_0_microseconds[5]\, Y => HIEFFPLA_NET_0_72132);
    
    HIEFFPLA_INST_0_65268 : AND2B
      port map(A => \Sensors_0_pressure_raw[6]\, B => 
        \Sensors_0_pressure_raw[12]\, Y => HIEFFPLA_NET_0_73430);
    
    HIEFFPLA_INST_0_59387 : MX2
      port map(A => HIEFFPLA_NET_0_74465, B => 
        HIEFFPLA_NET_0_74393, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74561);
    
    HIEFFPLA_INST_0_59595 : MX2
      port map(A => HIEFFPLA_NET_0_74419, B => 
        HIEFFPLA_NET_0_74412, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74533);
    
    \FMC_DA_pad[5]/U0/U1\ : IOTRI_OB_EB
      port map(D => \FMC_DA_c[5]\, E => \VCC\, DOUT => 
        \FMC_DA_pad[5]/U0/NET1\, EOUT => \FMC_DA_pad[5]/U0/NET2\);
    
    HIEFFPLA_INST_0_61270 : AX1
      port map(A => HIEFFPLA_NET_0_74244, B => 
        HIEFFPLA_NET_0_74250, C => 
        \General_Controller_0/state_seconds[16]_net_1\, Y => 
        HIEFFPLA_NET_0_74231);
    
    HIEFFPLA_INST_0_62986 : AO1A
      port map(A => HIEFFPLA_NET_0_73830, B => 
        HIEFFPLA_NET_0_74026, C => HIEFFPLA_NET_0_73851, Y => 
        HIEFFPLA_NET_0_73852);
    
    HIEFFPLA_INST_0_68211 : OR3A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\, B => 
        HIEFFPLA_NET_0_72703, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, Y => 
        HIEFFPLA_NET_0_72705);
    
    \General_Controller_0/state_seconds[18]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74229, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[18]_net_1\);
    
    \Communications_0/UART_0/rx_count[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75560, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75555, Q => 
        \Communications_0/UART_0/rx_count[1]_net_1\);
    
    HIEFFPLA_INST_0_69375 : XA1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[3]_net_1\, 
        B => HIEFFPLA_NET_0_72411, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72405);
    
    HIEFFPLA_INST_0_61985 : NAND2
      port map(A => \General_Controller_0/uc_rx_byte[3]_net_1\, B
         => \General_Controller_0/uc_rx_byte[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74082);
    
    HIEFFPLA_INST_0_68303 : XA1C
      port map(A => HIEFFPLA_NET_0_72690, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[3]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_72685);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/i2c_addr_1[1]\ : 
        DFN1E0
      port map(D => HIEFFPLA_NET_0_72994, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72774, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[1]\);
    
    \Timekeeper_0/milliseconds[23]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72101, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[23]\);
    
    HIEFFPLA_INST_0_70231 : AOI1C
      port map(A => HIEFFPLA_NET_0_72178, B => 
        HIEFFPLA_NET_0_72177, C => HIEFFPLA_NET_0_72273, Y => 
        HIEFFPLA_NET_0_72190);
    
    AFLSDF_INV_10 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_10\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/data_out_1[4]\ : 
        DFN1E1
      port map(D => HIEFFPLA_NET_0_73004, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72795, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[4]\);
    
    HIEFFPLA_INST_0_70673 : XOR2
      port map(A => \Timing_0/s_time[0]_net_1\, B => 
        HIEFFPLA_NET_0_72058, Y => HIEFFPLA_NET_0_72048);
    
    HIEFFPLA_INST_0_69316 : XA1B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        B => HIEFFPLA_NET_0_72380, C => HIEFFPLA_NET_0_72415, Y
         => HIEFFPLA_NET_0_72420);
    
    HIEFFPLA_INST_0_64181 : NOR3A
      port map(A => HIEFFPLA_NET_0_73751, B => 
        \General_Controller_0/uc_tx_state[12]_net_1\, C => 
        \General_Controller_0/uc_tx_state[14]_net_1\, Y => 
        HIEFFPLA_NET_0_73655);
    
    HIEFFPLA_INST_0_55468 : NOR2A
      port map(A => HIEFFPLA_NET_0_75497, B => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_75504);
    
    HIEFFPLA_INST_0_63052 : AXOI5
      port map(A => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_byte[4]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73840);
    
    \General_Controller_0/unit_id[6]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73990, Q => 
        \General_Controller_0_unit_id[6]\);
    
    \General_Controller_0/uc_send[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73769, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73601, Q => 
        \General_Controller_0_uc_send[0]\);
    
    HIEFFPLA_INST_0_70094 : AO1B
      port map(A => \Eject_Signal_Debounce_0/old_1kHz_i_0\, B => 
        \m_time[7]\, C => HIEFFPLA_NET_0_72236, Y => 
        HIEFFPLA_NET_0_72221);
    
    HIEFFPLA_INST_0_55519 : AND2
      port map(A => HIEFFPLA_NET_0_75488, B => 
        HIEFFPLA_NET_0_75453, Y => HIEFFPLA_NET_0_75489);
    
    HIEFFPLA_INST_0_55082 : NOR3A
      port map(A => \Communications_0/UART_0/rx_state[1]_net_1\, 
        B => \Communications_0/UART_0/rx_clk_count[25]_net_1\, C
         => \Communications_0/UART_0/rx_clk_count[26]_net_1\, Y
         => HIEFFPLA_NET_0_75595);
    
    \GS_Readout_0/state[6]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74599, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/state[6]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[3]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[3]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[3]\);
    
    HIEFFPLA_INST_0_55496 : NOR3A
      port map(A => GS_Readout_0_wen, B => 
        \Communications_0/UART_0/tx_state[0]_net_1\, C => 
        \Communications_0/UART_0/tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75497);
    
    \FPGA_BUF_INT_pad/U0/U0\ : IOPAD_TRI
      port map(D => \FPGA_BUF_INT_pad/U0/NET1\, E => 
        \FPGA_BUF_INT_pad/U0/NET2\, PAD => FPGA_BUF_INT);
    
    HIEFFPLA_INST_0_61228 : OR3B
      port map(A => HIEFFPLA_NET_0_74250, B => 
        \General_Controller_0/state_seconds[16]_net_1\, C => 
        HIEFFPLA_NET_0_74244, Y => HIEFFPLA_NET_0_74243);
    
    \General_Controller_0/state_seconds[11]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74238, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[11]_net_1\);
    
    HIEFFPLA_INST_0_67791 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        B => HIEFFPLA_NET_0_72765, C => HIEFFPLA_NET_0_72900, Y
         => HIEFFPLA_NET_0_72801);
    
    HIEFFPLA_INST_0_63031 : AO1
      port map(A => HIEFFPLA_NET_0_73825, B => 
        HIEFFPLA_NET_0_73783, C => HIEFFPLA_NET_0_73945, Y => 
        HIEFFPLA_NET_0_73844);
    
    HIEFFPLA_INST_0_66616 : AND3
      port map(A => HIEFFPLA_NET_0_73107, B => 
        HIEFFPLA_NET_0_73038, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[7]\, 
        Y => HIEFFPLA_NET_0_73082);
    
    HIEFFPLA_INST_0_66145 : MX2
      port map(A => \Science_0/DAC_SET_0/vector[16]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73196);
    
    HIEFFPLA_INST_0_69353 : NAND2B
      port map(A => HIEFFPLA_NET_0_72411, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72410);
    
    HIEFFPLA_INST_0_66779 : NOR3A
      port map(A => HIEFFPLA_NET_0_73044, B => 
        HIEFFPLA_NET_0_73027, C => HIEFFPLA_NET_0_73024, Y => 
        HIEFFPLA_NET_0_73036);
    
    HIEFFPLA_INST_0_67703 : AND3C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        B => HIEFFPLA_NET_0_72944, C => HIEFFPLA_NET_0_72942, Y
         => HIEFFPLA_NET_0_72819);
    
    \Science_0/ADC_READ_0/state[6]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_73237, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => \Science_0/ADC_READ_0/countere\);
    
    \Science_0/ADC_READ_0/data_a[16]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[16]_net_1\);
    
    HIEFFPLA_INST_0_55205 : OA1A
      port map(A => HIEFFPLA_NET_0_75558, B => 
        HIEFFPLA_NET_0_75564, C => 
        \Communications_0/UART_0/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75560);
    
    HIEFFPLA_INST_0_58149 : AO1
      port map(A => \Sensors_0_mag_time[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75146, Y => HIEFFPLA_NET_0_74839);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]\ : 
        DFN1P1
      port map(D => HIEFFPLA_NET_0_72746, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\);
    
    HIEFFPLA_INST_0_57059 : AOI1C
      port map(A => HIEFFPLA_NET_0_74887, B => 
        HIEFFPLA_NET_0_75032, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75174);
    
    HIEFFPLA_INST_0_65015 : OR2A
      port map(A => HIEFFPLA_NET_0_73482, B => 
        HIEFFPLA_NET_0_73487, Y => HIEFFPLA_NET_0_73488);
    
    HIEFFPLA_INST_0_67058 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[3]\, 
        B => \Sensors_0/Accelerometer_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72975);
    
    HIEFFPLA_INST_0_64614 : OR3A
      port map(A => HIEFFPLA_NET_0_73596, B => 
        \General_Controller_0/uc_tx_state[0]_net_1\, C => 
        \General_Controller_0/uc_tx_state[14]_net_1\, Y => 
        HIEFFPLA_NET_0_73586);
    
    \Communications_0/UART_0/tx_clk_count[7]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75519, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_clk_count_i_0[7]\);
    
    HIEFFPLA_INST_0_58605 : AND2B
      port map(A => \GS_Readout_0/prevState[0]_net_1\, B => 
        \GS_Readout_0/prevState[7]_net_1\, Y => 
        HIEFFPLA_NET_0_74723);
    
    HIEFFPLA_INST_0_55671 : OA1A
      port map(A => HIEFFPLA_NET_0_75447, B => 
        HIEFFPLA_NET_0_75453, C => 
        \Communications_0/UART_1/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75449);
    
    HIEFFPLA_INST_0_69030 : NAND2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        B => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72491);
    
    HIEFFPLA_INST_0_60916 : NOR3B
      port map(A => HIEFFPLA_NET_0_74028, B => 
        HIEFFPLA_NET_0_74325, C => HIEFFPLA_NET_0_74323, Y => 
        HIEFFPLA_NET_0_74320);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_0[11]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74772, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\);
    
    HIEFFPLA_INST_0_69058 : AOI1D
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[6]_net_1\, 
        C => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, Y => 
        HIEFFPLA_NET_0_72483);
    
    HIEFFPLA_INST_0_62413 : XNOR2
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73987);
    
    HIEFFPLA_INST_0_66170 : NOR2A
      port map(A => \Science_0/DAC_SET_0/vector[6]_net_1\, B => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73189);
    
    HIEFFPLA_INST_0_66882 : XOR2
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        B => HIEFFPLA_NET_0_73054, Y => HIEFFPLA_NET_0_73011);
    
    HIEFFPLA_INST_0_64912 : MX2
      port map(A => HIEFFPLA_NET_0_73507, B => FRAM_SDA_in, S => 
        \I2C_PassThrough_0.state[2]\, Y => HIEFFPLA_NET_0_73512);
    
    HIEFFPLA_INST_0_61331 : OR3B
      port map(A => 
        \General_Controller_0/state_seconds[18]_net_1\, B => 
        \General_Controller_0/state_seconds[17]_net_1\, C => 
        HIEFFPLA_NET_0_74243, Y => HIEFFPLA_NET_0_74215);
    
    HIEFFPLA_INST_0_69747 : NOR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        B => \Sensors_0/Pressure_Sensor_0/state[8]\, C => 
        HIEFFPLA_NET_0_72285, Y => HIEFFPLA_NET_0_72317);
    
    \Science_0/DAC_SET_0/cnt[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73219, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/cnt[0]_net_1\);
    
    HIEFFPLA_INST_0_70653 : XA1B
      port map(A => \Timing_0/s_count[4]_net_1\, B => 
        HIEFFPLA_NET_0_72021, C => HIEFFPLA_NET_0_72058, Y => 
        HIEFFPLA_NET_0_72053);
    
    HIEFFPLA_INST_0_58294 : AO1
      port map(A => \Science_0_exp_packet_0[41]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_75087, Y => HIEFFPLA_NET_0_74809);
    
    \Science_0/SET_LP_GAIN_0/state[4]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73155, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/state[4]_net_1\);
    
    HIEFFPLA_INST_0_67072 : NAND2B
      port map(A => HIEFFPLA_NET_0_72970, B => 
        HIEFFPLA_NET_0_72741, Y => HIEFFPLA_NET_0_72971);
    
    HIEFFPLA_INST_0_61726 : AOI1B
      port map(A => 
        \General_Controller_0/sweep_table_read_wait[30]_net_1\, B
         => 
        \General_Controller_0/sweep_table_read_wait[31]_net_1\, C
         => HIEFFPLA_NET_0_73779, Y => HIEFFPLA_NET_0_74153);
    
    \Timekeeper_0/milliseconds[15]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72110, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[15]\);
    
    HIEFFPLA_INST_0_57678 : AOI1
      port map(A => \Science_0_exp_packet_0[49]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74824, Y => HIEFFPLA_NET_0_74973);
    
    HIEFFPLA_INST_0_70037 : NOR2A
      port map(A => HIEFFPLA_NET_0_72301, B => 
        HIEFFPLA_NET_0_72235, Y => HIEFFPLA_NET_0_72238);
    
    \Science_0/ADC_READ_0/exp_packet_1[25]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[9]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[25]\);
    
    HIEFFPLA_INST_0_58975 : OA1A
      port map(A => HIEFFPLA_NET_0_74517, B => 
        HIEFFPLA_NET_0_74426, C => \GS_Readout_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_74645);
    
    HIEFFPLA_INST_0_56796 : MX2
      port map(A => HIEFFPLA_NET_0_75172, B => 
        HIEFFPLA_NET_0_75028, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75209);
    
    \Timekeeper_0/microseconds[8]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72129, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[8]\);
    
    HIEFFPLA_INST_0_61782 : XOR2
      port map(A => HIEFFPLA_NET_0_74148, B => 
        \General_Controller_0/sweep_table_sweep_cnt[3]_net_1\, Y
         => HIEFFPLA_NET_0_74135);
    
    HIEFFPLA_INST_0_55091 : NOR3A
      port map(A => HIEFFPLA_NET_0_75584, B => 
        \Communications_0/UART_0/rx_state[0]_net_1\, C => 
        \Communications_0/UART_0/rx_clk_count[23]_net_1\, Y => 
        HIEFFPLA_NET_0_75593);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/temp[4]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72907, Q => 
        \Sensors_0_acc_temp[4]\);
    
    \General_Controller_0/sweep_table_probe_id[7]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73924, Q => 
        \General_Controller_0/sweep_table_probe_id[7]_net_1\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/s_ack_error\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_73048, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73102, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\);
    
    HIEFFPLA_INST_0_58577 : AX1
      port map(A => HIEFFPLA_NET_0_74726, B => 
        \Eject_Signal_Debounce_0/ms_cnt[2]_net_1\, C => 
        \Eject_Signal_Debounce_0/ms_cnt[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74731);
    
    HIEFFPLA_INST_0_60680 : AND3
      port map(A => HIEFFPLA_NET_0_74341, B => 
        HIEFFPLA_NET_0_74342, C => HIEFFPLA_NET_0_74531, Y => 
        HIEFFPLA_NET_0_74377);
    
    \General_Controller_0/uc_rx_prev_state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74057, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_prev_state[1]_net_1\);
    
    HIEFFPLA_INST_0_70648 : XA1B
      port map(A => HIEFFPLA_NET_0_72025, B => 
        \Timing_0/s_count[3]_net_1\, C => HIEFFPLA_NET_0_72058, Y
         => HIEFFPLA_NET_0_72054);
    
    HIEFFPLA_INST_0_68386 : NAND3B
      port map(A => HIEFFPLA_NET_0_72647, B => 
        HIEFFPLA_NET_0_72651, C => HIEFFPLA_NET_0_72660, Y => 
        HIEFFPLA_NET_0_72661);
    
    HIEFFPLA_INST_0_60763 : MX2
      port map(A => HIEFFPLA_NET_0_74516, B => 
        HIEFFPLA_NET_0_74378, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74362);
    
    HIEFFPLA_INST_0_70111 : AOI1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\, 
        C => HIEFFPLA_NET_0_72271, Y => HIEFFPLA_NET_0_72216);
    
    HIEFFPLA_INST_0_58847 : AO1
      port map(A => HIEFFPLA_NET_0_74633, B => 
        HIEFFPLA_NET_0_74574, C => HIEFFPLA_NET_0_74669, Y => 
        HIEFFPLA_NET_0_74674);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[8]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[8]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[8]\);
    
    HIEFFPLA_INST_0_57140 : AND2
      port map(A => \Sensors_0_pressure_temp_raw[20]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75157);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[19]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[19]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[19]\);
    
    \Science_0/ADC_READ_0/cnt1up[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73391, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1up[4]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/data_out[28]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75215, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[28]\);
    
    HIEFFPLA_INST_0_62944 : NAND3C
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73861);
    
    HIEFFPLA_INST_0_70768 : AO1
      port map(A => HIEFFPLA_NET_0_72200, B => 
        HIEFFPLA_NET_0_72230, C => HIEFFPLA_NET_0_72201, Y => 
        HIEFFPLA_NET_0_72016);
    
    HIEFFPLA_INST_0_59643 : MX2
      port map(A => HIEFFPLA_NET_0_74555, B => 
        HIEFFPLA_NET_0_74501, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74527);
    
    HIEFFPLA_INST_0_63081 : AOI1D
      port map(A => HIEFFPLA_NET_0_73888, B => 
        HIEFFPLA_NET_0_73831, C => HIEFFPLA_NET_0_73780, Y => 
        HIEFFPLA_NET_0_73833);
    
    HIEFFPLA_INST_0_63036 : AND3
      port map(A => HIEFFPLA_NET_0_73775, B => 
        HIEFFPLA_NET_0_74070, C => HIEFFPLA_NET_0_73956, Y => 
        HIEFFPLA_NET_0_73843);
    
    HIEFFPLA_INST_0_55939 : AND3
      port map(A => \Communications_0/UART_1/tx_count[0]_net_1\, 
        B => \Communications_0/UART_1/tx_count[1]_net_1\, C => 
        \Communications_0/UART_1/tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75390);
    
    HIEFFPLA_INST_0_56311 : AO13
      port map(A => HIEFFPLA_NET_0_75339, B => 
        HIEFFPLA_NET_0_75312, C => HIEFFPLA_NET_0_75274, Y => 
        HIEFFPLA_NET_0_75311);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_WADDR[4]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75315, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\);
    
    HIEFFPLA_INST_0_57447 : AO1
      port map(A => \Sensors_0_acc_z[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74866, Y => HIEFFPLA_NET_0_75043);
    
    HIEFFPLA_INST_0_56897 : MX2
      port map(A => HIEFFPLA_NET_0_74993, B => 
        HIEFFPLA_NET_0_74921, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75198);
    
    \GS_Readout_0/prevState[7]\ : DFN1E0P1
      port map(D => \GS_Readout_0/state[7]_net_1\, CLK => 
        CLKINT_0_Y_0, PRE => CLKINT_1_Y, E => 
        \GS_Readout_0/state[6]_net_1\, Q => 
        \GS_Readout_0/prevState[7]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/data_out[31]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75211, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[31]\);
    
    HIEFFPLA_INST_0_68752 : NAND3C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, Y
         => HIEFFPLA_NET_0_72570);
    
    HIEFFPLA_INST_0_68568 : AO1
      port map(A => HIEFFPLA_NET_0_72584, B => 
        HIEFFPLA_NET_0_72663, C => HIEFFPLA_NET_0_72614, Y => 
        HIEFFPLA_NET_0_72615);
    
    \Science_0/ADC_READ_0/state[1]\ : DFN1C1
      port map(D => \Science_0/ADC_READ_0/state[2]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => 
        \Science_0/ADC_READ_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_59545 : MX2
      port map(A => \Science_0_chan6_data[7]\, B => 
        \Science_0_chan6_data[11]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74540);
    
    HIEFFPLA_INST_0_58038 : AND2
      port map(A => \Sensors_0_gyro_x[14]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_74871);
    
    \General_Controller_0/uc_rx_substate[0]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_73774, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_substate[0]_net_1\);
    
    HIEFFPLA_INST_0_57143 : AND2
      port map(A => \Sensors_0_pressure_temp_raw[23]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75155);
    
    HIEFFPLA_INST_0_59663 : MX2
      port map(A => HIEFFPLA_NET_0_74399, B => 
        HIEFFPLA_NET_0_74425, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74525);
    
    HIEFFPLA_INST_0_58254 : AO1
      port map(A => \Sensors_0_gyro_time[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75111, Y => HIEFFPLA_NET_0_74819);
    
    \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[0]\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72688, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72618, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[0]_net_1\);
    
    HIEFFPLA_INST_0_62781 : NOR2A
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73905);
    
    HIEFFPLA_INST_0_62678 : AO1A
      port map(A => \General_Controller_0/uc_rx_state[1]_net_1\, 
        B => HIEFFPLA_NET_0_73796, C => HIEFFPLA_NET_0_74020, Y
         => HIEFFPLA_NET_0_73930);
    
    HIEFFPLA_INST_0_57821 : AOI1C
      port map(A => HIEFFPLA_NET_0_74768, B => 
        HIEFFPLA_NET_0_75165, C => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        Y => HIEFFPLA_NET_0_74934);
    
    HIEFFPLA_INST_0_70435 : AX1C
      port map(A => \Timekeeper_0_microseconds[5]\, B => 
        HIEFFPLA_NET_0_72156, C => \Timekeeper_0_microseconds[6]\, 
        Y => HIEFFPLA_NET_0_72131);
    
    HIEFFPLA_INST_0_60391 : MX2
      port map(A => \Science_0_chan5_data[3]\, B => 
        \Science_0_chan5_data[7]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74422);
    
    HIEFFPLA_INST_0_57883 : AO1
      port map(A => \Science_0_exp_packet_0[79]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75135, Y => HIEFFPLA_NET_0_74916);
    
    HIEFFPLA_INST_0_66315 : AND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73148);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[0]\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72300, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72221, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[0]_net_1\);
    
    \General_Controller_0/sweep_table_points[10]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[10]_net_1\);
    
    \CLOCK_pad/U0/U0\ : IOPAD_IN
      port map(PAD => CLOCK, Y => \CLOCK_pad/U0/NET1\);
    
    \Science_0/ADC_READ_0/cnt4dn[7]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73311, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4dn[7]_net_1\);
    
    \LDSDI_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => LDSDI_c, E => \VCC\, DOUT => 
        \LDSDI_pad/U0/NET1\, EOUT => \LDSDI_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_57703 : AO1
      port map(A => \Sensors_0_pressure_raw[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74846, Y => HIEFFPLA_NET_0_74965);
    
    HIEFFPLA_INST_0_71215 : OA1C
      port map(A => \Communications_0/UART_0_rx_rdy\, B => 
        \Communications_0/FFU_Command_Checker_0/state[1]_net_1\, 
        C => HIEFFPLA_NET_0_71971, Y => HIEFFPLA_NET_0_75622);
    
    HIEFFPLA_INST_0_69419 : AO1A
      port map(A => PRESSURE_SCL_c, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        C => HIEFFPLA_NET_0_72341, Y => HIEFFPLA_NET_0_72393);
    
    HIEFFPLA_INST_0_63908 : MX2
      port map(A => HIEFFPLA_NET_0_73668, B => 
        HIEFFPLA_NET_0_73661, S => HIEFFPLA_NET_0_73594, Y => 
        HIEFFPLA_NET_0_73691);
    
    HIEFFPLA_INST_0_62204 : AND2
      port map(A => HIEFFPLA_NET_0_73943, B => 
        Communications_0_uc_rx_rdy, Y => HIEFFPLA_NET_0_74030);
    
    HIEFFPLA_INST_0_69610 : NOR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[2]_net_1\, 
        B => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72350);
    
    HIEFFPLA_INST_0_55447 : NOR3B
      port map(A => \Communications_0/UART_0/tx_count[2]_net_1\, 
        B => \Communications_0/UART_0/tx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_75528, Y => HIEFFPLA_NET_0_75510);
    
    HIEFFPLA_INST_0_59737 : MX2
      port map(A => \Sensors_0_pressure_temp_raw[13]\, B => 
        \Sensors_0_pressure_temp_raw[17]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74515);
    
    HIEFFPLA_INST_0_56622 : MX2
      port map(A => HIEFFPLA_NET_0_75198, B => 
        HIEFFPLA_NET_0_75067, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75231);
    
    HIEFFPLA_INST_0_55053 : NOR3A
      port map(A => \Communications_0/UART_0/rx_count[0]_net_1\, 
        B => \Communications_0/UART_0/rx_count[2]_net_1\, C => 
        \Communications_0/UART_0/rx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75602);
    
    HIEFFPLA_INST_0_67900 : AND3C
      port map(A => HIEFFPLA_NET_0_72757, B => 
        HIEFFPLA_NET_0_72775, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72777);
    
    HIEFFPLA_INST_0_59056 : AND3
      port map(A => HIEFFPLA_NET_0_74481, B => 
        HIEFFPLA_NET_0_74459, C => HIEFFPLA_NET_0_74619, Y => 
        HIEFFPLA_NET_0_74624);
    
    \Science_0/ADC_READ_0/exp_packet_1[11]\ : DFN1E0
      port map(D => \AFLSDF_INV_13\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[11]\);
    
    HIEFFPLA_INST_0_66107 : AO1A
      port map(A => \Science_0/DAC_SET_0/state[3]_net_1\, B => 
        HIEFFPLA_NET_0_73206, C => HIEFFPLA_NET_0_73205, Y => 
        HIEFFPLA_NET_0_73208);
    
    HIEFFPLA_INST_0_65622 : AND2
      port map(A => HIEFFPLA_NET_0_73322, B => 
        \Science_0/ADC_READ_0/cnt4dn[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73327);
    
    HIEFFPLA_INST_0_62353 : AOI1C
      port map(A => HIEFFPLA_NET_0_73776, B => 
        HIEFFPLA_NET_0_74019, C => HIEFFPLA_NET_0_73998, Y => 
        HIEFFPLA_NET_0_73999);
    
    HIEFFPLA_INST_0_57893 : AO1
      port map(A => \Science_0_exp_packet_0[64]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75134, Y => HIEFFPLA_NET_0_74913);
    
    HIEFFPLA_INST_0_70706 : NAND3
      port map(A => HIEFFPLA_NET_0_72035, B => 
        \Timing_0/s_time[7]_net_1\, C => 
        \Timing_0/s_time[4]_net_1\, Y => HIEFFPLA_NET_0_72036);
    
    HIEFFPLA_INST_0_60728 : NOR2A
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74368);
    
    HIEFFPLA_INST_0_59377 : MX2
      port map(A => HIEFFPLA_NET_0_74424, B => 
        HIEFFPLA_NET_0_74447, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74562);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[6]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72463, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[6]_net_1\);
    
    \General_Controller_0/sweep_table_samples_per_point[14]\ : 
        DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[14]_net_1\);
    
    HIEFFPLA_INST_0_57637 : AO1
      port map(A => \Sensors_0_pressure_raw[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74794, Y => HIEFFPLA_NET_0_74985);
    
    AFLSDF_INV_29 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_29\);
    
    HIEFFPLA_INST_0_56837 : MX2
      port map(A => HIEFFPLA_NET_0_75167, B => 
        HIEFFPLA_NET_0_75016, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75205);
    
    HIEFFPLA_INST_0_57749 : AO1
      port map(A => \Sensors_0_pressure_raw[18]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, C
         => HIEFFPLA_NET_0_74953, Y => HIEFFPLA_NET_0_74954);
    
    \Data_Saving_0/Packet_Saver_0/data_out[23]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75221, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[23]\);
    
    \Communications_0/UART_1/tx_clk_count[3]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75408, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_clk_count_i_0[3]\);
    
    \Science_0/ADC_READ_0/chan3_data[8]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[8]\);
    
    HIEFFPLA_INST_0_56105 : XA1B
      port map(A => HIEFFPLA_NET_0_75366, B => 
        HIEFFPLA_NET_0_89701, C => HIEFFPLA_NET_0_89700, Y => 
        HIEFFPLA_NET_0_75346);
    
    HIEFFPLA_INST_0_58074 : AO1
      port map(A => \Sensors_0_gyro_y[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75156, Y => HIEFFPLA_NET_0_74863);
    
    HIEFFPLA_INST_0_55995 : XOR2
      port map(A => HIEFFPLA_NET_0_75321, B => 
        HIEFFPLA_NET_0_75288, Y => HIEFFPLA_NET_0_75374);
    
    \Science_0/ADC_READ_0/chan6_data[5]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[5]\);
    
    \Science_0/ADC_READ_0/chan0_data[5]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[5]\);
    
    HIEFFPLA_INST_0_63064 : AND3
      port map(A => HIEFFPLA_NET_0_73832, B => 
        HIEFFPLA_NET_0_73908, C => HIEFFPLA_NET_0_73907, Y => 
        HIEFFPLA_NET_0_73837);
    
    HIEFFPLA_INST_0_63692 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[2]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_nof_steps[2]_net_1\, S
         => \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73727);
    
    HIEFFPLA_INST_0_61278 : XA1C
      port map(A => 
        \General_Controller_0/state_seconds[18]_net_1\, B => 
        HIEFFPLA_NET_0_74255, C => HIEFFPLA_NET_0_74217, Y => 
        HIEFFPLA_NET_0_74229);
    
    HIEFFPLA_INST_0_69825 : NOR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[4]_net_1\, 
        B => HIEFFPLA_NET_0_72303, Y => HIEFFPLA_NET_0_72294);
    
    HIEFFPLA_INST_0_66808 : AO1
      port map(A => HIEFFPLA_NET_0_73101, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_73030);
    
    HIEFFPLA_INST_0_58865 : NOR3B
      port map(A => HIEFFPLA_NET_0_74496, B => 
        HIEFFPLA_NET_0_74617, C => HIEFFPLA_NET_0_74459, Y => 
        HIEFFPLA_NET_0_74670);
    
    HIEFFPLA_INST_0_68833 : AND3
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, C => 
        HIEFFPLA_NET_0_72545, Y => HIEFFPLA_NET_0_72546);
    
    \Data_Saving_0/Packet_Saver_0/data_out[16]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75229, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[16]\);
    
    HIEFFPLA_INST_0_68709 : NAND3C
      port map(A => HIEFFPLA_NET_0_72631, B => 
        HIEFFPLA_NET_0_72689, C => GYRO_SCL_c, Y => 
        HIEFFPLA_NET_0_72581);
    
    HIEFFPLA_INST_0_62058 : NOR3B
      port map(A => HIEFFPLA_NET_0_74038, B => 
        HIEFFPLA_NET_0_74060, C => HIEFFPLA_NET_0_74024, Y => 
        HIEFFPLA_NET_0_74061);
    
    \Science_0/ADC_READ_0/cnt2up[1]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73363, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2up[1]_net_1\);
    
    HIEFFPLA_INST_0_61476 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[52]\, B => 
        \Timekeeper_0_milliseconds[12]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74194);
    
    HIEFFPLA_INST_0_58775 : NOR3B
      port map(A => HIEFFPLA_NET_0_74552, B => 
        \GS_Readout_0/state[3]_net_1\, C => HIEFFPLA_NET_0_74474, 
        Y => HIEFFPLA_NET_0_74688);
    
    HIEFFPLA_INST_0_60513 : MX2
      port map(A => \Science_0_chan7_data[9]\, B => 
        \Science_0_chan6_data[1]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74403);
    
    HIEFFPLA_INST_0_60727 : NAND2B
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74369);
    
    \GS_Readout_0/state[7]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_74598, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => \GS_Readout_0/state[7]_net_1\);
    
    AFLSDF_INV_27 : INV
      port map(A => 
        \Communications_0/FFU_Command_Checker_0/state[0]_net_1\, 
        Y => \AFLSDF_INV_27\);
    
    HIEFFPLA_INST_0_59830 : MX2
      port map(A => HIEFFPLA_NET_0_74489, B => 
        HIEFFPLA_NET_0_74543, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74501);
    
    \Science_0/ADC_READ_0/cnt_chan[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73278, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/ADC_READ_0/cnt_chan[1]_net_1\);
    
    HIEFFPLA_INST_0_56524 : AND3
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[3]_net_1\, B
         => HIEFFPLA_NET_0_75256, C => 
        \Data_Saving_0/Interrupt_Generator_0/counter[4]_net_1\, Y
         => HIEFFPLA_NET_0_75254);
    
    HIEFFPLA_INST_0_60400 : MX2
      port map(A => HIEFFPLA_NET_0_74467, B => 
        HIEFFPLA_NET_0_74485, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74420);
    
    HIEFFPLA_INST_0_60711 : NOR2A
      port map(A => HIEFFPLA_NET_0_74527, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74372);
    
    HIEFFPLA_INST_0_61717 : MX2
      port map(A => \SweepTable_0_RD[9]\, B => 
        \SweepTable_1_RD[9]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74155);
    
    HIEFFPLA_INST_0_61201 : OR3B
      port map(A => 
        \General_Controller_0/state_seconds[10]_net_1\, B => 
        \General_Controller_0/state_seconds[11]_net_1\, C => 
        HIEFFPLA_NET_0_74241, Y => HIEFFPLA_NET_0_74251);
    
    HIEFFPLA_INST_0_64201 : NOR3A
      port map(A => HIEFFPLA_NET_0_73746, B => 
        \General_Controller_0/uc_tx_state[12]_net_1\, C => 
        \General_Controller_0/uc_tx_state[14]_net_1\, Y => 
        HIEFFPLA_NET_0_73650);
    
    \General_Controller_0/sweep_table_read_wait[31]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74151, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/sweep_table_read_wait[31]_net_1\);
    
    HIEFFPLA_INST_0_70532 : NOR2A
      port map(A => \s_clks_net_0[4]\, B => 
        \Timekeeper_0/old_1MHz_net_1\, Y => HIEFFPLA_NET_0_72092);
    
    HIEFFPLA_INST_0_66169 : NOR2A
      port map(A => \Science_0/DAC_SET_0/vector[5]_net_1\, B => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73190);
    
    \FRAM_SDA_pad/U0/U0\ : IOPAD_BI
      port map(D => \FRAM_SDA_pad/U0/NET1\, E => 
        \FRAM_SDA_pad/U0/NET2\, Y => \FRAM_SDA_pad/U0/NET3\, PAD
         => FRAM_SDA);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[16]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72280, Q => \Sensors_0_pressure_raw[16]\);
    
    \Science_0/ADC_READ_0/cnt1up[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73397, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1up[0]_net_1\);
    
    HIEFFPLA_INST_0_68085 : OR3A
      port map(A => HIEFFPLA_NET_0_72731, B => 
        HIEFFPLA_NET_0_72910, C => HIEFFPLA_NET_0_72732, Y => 
        HIEFFPLA_NET_0_72733);
    
    HIEFFPLA_INST_0_57264 : AND2
      port map(A => \Sensors_0_gyro_y[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75105);
    
    HIEFFPLA_INST_0_55443 : NAND2
      port map(A => \Communications_0/UART_0/tx_count[0]_net_1\, 
        B => \Communications_0/UART_0/tx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75511);
    
    \General_Controller_0/uc_send[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73767, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73601, Q => 
        \General_Controller_0_uc_send[2]\);
    
    HIEFFPLA_INST_0_66225 : MX2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G2[0]_net_1\, B
         => \Science_0/ADC_READ_0_G2[0]\, S => 
        \Science_0/SET_LP_GAIN_0/state[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73173);
    
    HIEFFPLA_INST_0_59022 : OR3A
      port map(A => \GS_Readout_0/state[5]_net_1\, B => 
        \GS_Readout_0/subState[0]_net_1\, C => 
        \GS_Readout_0/subState[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74634);
    
    \Science_0/ADC_READ_0/chan5_data[4]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[4]\);
    
    \AB_pad/U0/U0\ : IOPAD_IN
      port map(PAD => AB, Y => \AB_pad/U0/NET1\);
    
    \Communications_0/FFU_Command_Checker_0/rmu_oen\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75624, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/FFU_Command_Checker_0_rmu_oen\);
    
    HIEFFPLA_INST_0_67334 : AOI1
      port map(A => HIEFFPLA_NET_0_72751, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        C => HIEFFPLA_NET_0_72933, Y => HIEFFPLA_NET_0_72905);
    
    HIEFFPLA_INST_0_67759 : NOR3B
      port map(A => HIEFFPLA_NET_0_72738, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        C => HIEFFPLA_NET_0_72874, Y => HIEFFPLA_NET_0_72808);
    
    \Science_0/ADC_READ_0/chan0_data[10]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[10]\);
    
    HIEFFPLA_INST_0_64992 : XA1
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[1]_net_1\, 
        B => HIEFFPLA_NET_0_73449, C => HIEFFPLA_NET_0_73490, Y
         => HIEFFPLA_NET_0_73494);
    
    \Data_Saving_0/Packet_Saver_0/data_out[10]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75235, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[10]\);
    
    \Science_0/ADC_READ_0/state[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73239, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/ADC_READ_0/state[2]_net_1\);
    
    HIEFFPLA_INST_0_65501 : XA1
      port map(A => HIEFFPLA_NET_0_73367, B => 
        \Science_0/ADC_READ_0/cnt2up[3]_net_1\, C => 
        HIEFFPLA_NET_0_73366, Y => HIEFFPLA_NET_0_73361);
    
    HIEFFPLA_INST_0_56238 : XOR3
      port map(A => HIEFFPLA_NET_0_75312, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[4]\\\\\, C => 
        HIEFFPLA_NET_0_75273, Y => HIEFFPLA_NET_0_75327);
    
    AFLSDF_INV_1 : INV
      port map(A => \Data_Saving_0/FPGA_Buffer_0/MEMRENEG\, Y => 
        \AFLSDF_INV_1\);
    
    \GS_Readout_0/send[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74715, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74630, Q => 
        \GS_Readout_0_send[2]\);
    
    HIEFFPLA_INST_0_69759 : AOI1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        B => \Sensors_0/Pressure_Sensor_0/state[8]\, C => 
        HIEFFPLA_NET_0_72224, Y => HIEFFPLA_NET_0_72314);
    
    HIEFFPLA_INST_0_70540 : XOR2
      port map(A => \Timing_0/f_time[3]_net_1\, B => 
        HIEFFPLA_NET_0_72090, Y => HIEFFPLA_NET_0_72087);
    
    HIEFFPLA_INST_0_59294 : MX2
      port map(A => \Science_0_chan7_data[10]\, B => 
        \Science_0_chan6_data[2]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74573);
    
    \General_Controller_0/uc_send[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73765, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73601, Q => 
        \General_Controller_0_uc_send[4]\);
    
    HIEFFPLA_INST_0_62832 : NAND2B
      port map(A => \General_Controller_0/uc_rx_state[4]_net_1\, 
        B => \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73889);
    
    HIEFFPLA_INST_0_61776 : AX1
      port map(A => HIEFFPLA_NET_0_74128, B => 
        \General_Controller_0/sweep_table_sweep_cnt[13]_net_1\, C
         => 
        \General_Controller_0/sweep_table_sweep_cnt[15]_net_1\, Y
         => HIEFFPLA_NET_0_74138);
    
    HIEFFPLA_INST_0_62776 : AND2B
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73908);
    
    HIEFFPLA_INST_0_65647 : NOR2A
      port map(A => HIEFFPLA_NET_0_73274, B => 
        \Science_0/ADC_READ_0/cnt4dn[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73318);
    
    HIEFFPLA_INST_0_65231 : AND3C
      port map(A => HIEFFPLA_NET_0_73467, B => 
        HIEFFPLA_NET_0_73459, C => HIEFFPLA_NET_0_73438, Y => 
        HIEFFPLA_NET_0_73439);
    
    HIEFFPLA_INST_0_63884 : AND2
      port map(A => HIEFFPLA_NET_0_73664, B => 
        HIEFFPLA_NET_0_73594, Y => HIEFFPLA_NET_0_73695);
    
    \Timekeeper_0/milliseconds[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72099, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[3]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[13]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72281, Q => \Sensors_0_pressure_raw[13]\);
    
    HIEFFPLA_INST_0_67150 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72951);
    
    \General_Controller_0/old_status_packet_clk\ : DFN1P1
      port map(D => \AFLSDF_INV_14\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => 
        \General_Controller_0/old_status_packet_clk_i_0\);
    
    HIEFFPLA_INST_0_68680 : AND2B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_i2c_repeat_start\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0/state[2]_net_1\, Y
         => HIEFFPLA_NET_0_72590);
    
    HIEFFPLA_INST_0_55970 : NOR3A
      port map(A => General_Controller_0_uc_wen, B => 
        \Communications_0/UART_1/tx_state[0]_net_1\, C => 
        \Communications_0/UART_1/tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75381);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73033, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\);
    
    HIEFFPLA_INST_0_57971 : AO1
      port map(A => \Science_0_exp_packet_0[25]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74787, Y => HIEFFPLA_NET_0_74890);
    
    HIEFFPLA_INST_0_69422 : AO1D
      port map(A => HIEFFPLA_NET_0_72388, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        C => HIEFFPLA_NET_0_72391, Y => HIEFFPLA_NET_0_72392);
    
    HIEFFPLA_INST_0_65621 : AO1
      port map(A => HIEFFPLA_NET_0_73321, B => 
        HIEFFPLA_NET_0_73325, C => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_73328);
    
    \Communications_0/UART_0/tx_clk_count[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75525, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_clk_count[1]_net_1\);
    
    HIEFFPLA_INST_0_62783 : NOR3A
      port map(A => HIEFFPLA_NET_0_73906, B => 
        \General_Controller_0/uc_rx_state[3]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73904);
    
    \Science_0/SET_LP_GAIN_0/state[7]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73152, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/state[7]_net_1\);
    
    HIEFFPLA_INST_0_66003 : NAND2B
      port map(A => \Science_0/ADC_READ_0/countere\, B => 
        HIEFFPLA_NET_0_73238, Y => HIEFFPLA_NET_0_73241);
    
    HIEFFPLA_INST_0_70676 : AX1C
      port map(A => HIEFFPLA_NET_0_72033, B => 
        \Timing_0/s_time[2]_net_1\, C => \s_clks_net_0[18]\, Y
         => HIEFFPLA_NET_0_72047);
    
    HIEFFPLA_INST_0_64975 : AND3C
      port map(A => HIEFFPLA_NET_0_73496, B => 
        \Pressure_Signal_Debounce_0/ms_cnt[1]_net_1\, C => 
        \Pressure_Signal_Debounce_0/ms_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73497);
    
    HIEFFPLA_INST_0_66090 : AO1
      port map(A => LDCLK_c, B => HIEFFPLA_NET_0_73222, C => 
        HIEFFPLA_NET_0_73226, Y => HIEFFPLA_NET_0_73211);
    
    HIEFFPLA_INST_0_58495 : OR3A
      port map(A => \Eject_Signal_Debounce_0/ms_cnt[1]_net_1\, B
         => HIEFFPLA_NET_0_74748, C => 
        \Eject_Signal_Debounce_0/ms_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74749);
    
    HIEFFPLA_INST_0_67990 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => HIEFFPLA_NET_0_72739, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72760);
    
    HIEFFPLA_INST_0_61540 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[60]\, B => 
        \Timekeeper_0_milliseconds[20]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74186);
    
    \Science_0/ADC_READ_0/chan2_data[2]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[2]\);
    
    HIEFFPLA_INST_0_63812 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[6]_net_1\, 
        B => \General_Controller_0/sweep_table_points[6]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73707);
    
    HIEFFPLA_INST_0_63456 : MX2
      port map(A => HIEFFPLA_NET_0_73686, B => 
        HIEFFPLA_NET_0_73678, S => HIEFFPLA_NET_0_73621, Y => 
        HIEFFPLA_NET_0_73761);
    
    \Science_0/DAC_SET_0/vector[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73189, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[7]_net_1\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/data_out[5]\ : DFN0E1C1
      port map(D => GYRO_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72677, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[5]\);
    
    HIEFFPLA_INST_0_68545 : MX2
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, B => 
        HIEFFPLA_NET_0_72623, S => GYRO_SCL_c, Y => 
        HIEFFPLA_NET_0_72621);
    
    HIEFFPLA_INST_0_68372 : NOR2A
      port map(A => HIEFFPLA_NET_0_72698, B => 
        HIEFFPLA_NET_0_72700, Y => HIEFFPLA_NET_0_72666);
    
    HIEFFPLA_INST_0_69788 : OR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[3]_net_1\, 
        B => HIEFFPLA_NET_0_72307, Y => HIEFFPLA_NET_0_72303);
    
    HIEFFPLA_INST_0_67678 : NOR3B
      port map(A => HIEFFPLA_NET_0_72743, B => 
        HIEFFPLA_NET_0_72821, C => HIEFFPLA_NET_0_72792, Y => 
        HIEFFPLA_NET_0_72825);
    
    HIEFFPLA_INST_0_62599 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => HIEFFPLA_NET_0_73889, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73948);
    
    HIEFFPLA_INST_0_55065 : AND2
      port map(A => \Communications_0/UART_0/rx_count[2]_net_1\, 
        B => \Communications_0/UART_0/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75599);
    
    HIEFFPLA_INST_0_66337 : NOR3B
      port map(A => HIEFFPLA_NET_0_73059, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[3]_net_1\, 
        C => HIEFFPLA_NET_0_73143, Y => HIEFFPLA_NET_0_73142);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[2]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72489, Q => 
        \Sensors_0_gyro_z[2]\);
    
    HIEFFPLA_INST_0_70614 : AX1C
      port map(A => \Timing_0/m_time[0]_net_1\, B => 
        HIEFFPLA_NET_0_72083, C => \Timing_0/m_time[1]_net_1\, Y
         => HIEFFPLA_NET_0_72064);
    
    \General_Controller_0/command[5]\ : DFN1E1
      port map(D => \Communications_0_ext_recv[5]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74300, Q => 
        \General_Controller_0/command[5]_net_1\);
    
    \Science_0/ADC_READ_0/cnt1up[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73396, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1up[1]_net_1\);
    
    HIEFFPLA_INST_0_60338 : MX2
      port map(A => \Science_0_chan5_data[9]\, B => 
        \Science_0_chan4_data[1]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74430);
    
    HIEFFPLA_INST_0_64645 : NOR3B
      port map(A => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, B => 
        HIEFFPLA_NET_0_74325, C => HIEFFPLA_NET_0_73552, Y => 
        HIEFFPLA_NET_0_73578);
    
    HIEFFPLA_INST_0_70153 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[5]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72207);
    
    \Science_0/ADC_READ_0/exp_packet_1[41]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[7]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[41]\);
    
    HIEFFPLA_INST_0_88368 : AO18
      port map(A => HIEFFPLA_NET_0_75304, B => 
        HIEFFPLA_NET_0_75320, C => HIEFFPLA_NET_0_75288, Y => 
        HIEFFPLA_NET_0_88385);
    
    \General_Controller_0/constant_bias_voltage_0[6]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[6]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[6]_net_1\);
    
    HIEFFPLA_INST_0_70972 : XA1B
      port map(A => \Science_0/ADC_READ_0/data_b[12]_net_1\, B
         => \Science_0/ADC_READ_0/data_b[15]_net_1\, C => 
        HIEFFPLA_NET_0_71997, Y => HIEFFPLA_NET_0_73275);
    
    HIEFFPLA_INST_0_69787 : OA1C
      port map(A => HIEFFPLA_NET_0_72302, B => 
        HIEFFPLA_NET_0_72311, C => HIEFFPLA_NET_0_72235, Y => 
        HIEFFPLA_NET_0_72304);
    
    \Science_0/ADC_READ_0/chan7_data[5]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[5]\);
    
    HIEFFPLA_INST_0_70882 : OA1C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, B
         => HIEFFPLA_NET_0_72876, C => HIEFFPLA_NET_0_72005, Y
         => HIEFFPLA_NET_0_72755);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[3]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72279, Q => 
        \Sensors_0_pressure_temp_raw[3]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[10]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[10]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[10]\);
    
    \Science_0/ADC_READ_0/cnt4dn[1]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73317, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4dn[1]_net_1\);
    
    HIEFFPLA_INST_0_70350 : AOI1D
      port map(A => General_Controller_0_st_ren1, B => 
        \SweepTable_0/WEBP\, C => 
        \General_Controller_0_st_raddr_1[7]\, Y => 
        \TableSelect_0_RADDR[7]\);
    
    \Timekeeper_0/microseconds[23]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72136, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[23]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/i2c_addr_1[0]\ : 
        DFN1E0
      port map(D => HIEFFPLA_NET_0_72996, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72774, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[0]\);
    
    HIEFFPLA_INST_0_57023 : AOI1C
      port map(A => HIEFFPLA_NET_0_74889, B => 
        HIEFFPLA_NET_0_75039, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75180);
    
    HIEFFPLA_INST_0_57542 : AOI1
      port map(A => \Science_0_exp_packet_0[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_75014, Y => HIEFFPLA_NET_0_75015);
    
    HIEFFPLA_INST_0_64091 : MX2
      port map(A => HIEFFPLA_NET_0_73635, B => 
        HIEFFPLA_NET_0_73627, S => HIEFFPLA_NET_0_73585, Y => 
        HIEFFPLA_NET_0_73672);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_2\ : DFN1C0
      port map(D => \VCC\, CLK => CLKINT_2_Y, CLR => 
        \AFLSDF_INV_15\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_2_Q\);
    
    HIEFFPLA_INST_0_69186 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        B => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, 
        C => HIEFFPLA_NET_0_72540, Y => HIEFFPLA_NET_0_72452);
    
    \Science_0/ADC_READ_0/cnt3dn[3]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73344, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3dn[3]_net_1\);
    
    \Science_0/ADC_READ_0/chan1_data[0]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[0]\);
    
    HIEFFPLA_INST_0_69612 : AND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[5]_net_1\, 
        B => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72348);
    
    \GS_Readout_0/send[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74712, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74630, Q => 
        \GS_Readout_0_send[5]\);
    
    HIEFFPLA_INST_0_70212 : AND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[4]_net_1\, 
        C => HIEFFPLA_NET_0_72240, Y => HIEFFPLA_NET_0_72194);
    
    HIEFFPLA_INST_0_68435 : AND2
      port map(A => HIEFFPLA_NET_0_72648, B => 
        \Sensors_0.Gyro_0.I2C_Master_0.sda_1\, Y => 
        HIEFFPLA_NET_0_72651);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRYSYNC[4]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_3_Q\, CLK
         => CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[4]\\\\\);
    
    HIEFFPLA_INST_0_62619 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[1]_net_1\, 
        B => HIEFFPLA_NET_0_73889, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73943);
    
    \Timekeeper_0/old_1MHz\ : DFN1E0
      port map(D => \s_clks_net_0[4]\, CLK => CLKINT_0_Y_0, E => 
        CLKINT_1_Y, Q => \Timekeeper_0/old_1MHz_net_1\);
    
    HIEFFPLA_INST_0_65611 : AX1C
      port map(A => \Science_0/ADC_READ_0/cnt3up[2]_net_1\, B => 
        HIEFFPLA_NET_0_73337, C => 
        \Science_0/ADC_READ_0/cnt3up[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73331);
    
    HIEFFPLA_INST_0_69161 : NAND3C
      port map(A => HIEFFPLA_NET_0_72446, B => 
        HIEFFPLA_NET_0_72443, C => HIEFFPLA_NET_0_72442, Y => 
        HIEFFPLA_NET_0_72457);
    
    HIEFFPLA_INST_0_66366 : AX1E
      port map(A => HIEFFPLA_NET_0_73010, B => 
        HIEFFPLA_NET_0_73054, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73137);
    
    HIEFFPLA_INST_0_68017 : NOR3A
      port map(A => HIEFFPLA_NET_0_72738, B => 
        HIEFFPLA_NET_0_72939, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72753);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[9]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[9]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[9]\);
    
    HIEFFPLA_INST_0_65029 : AO1B
      port map(A => HIEFFPLA_NET_0_73446, B => 
        HIEFFPLA_NET_0_73477, C => HIEFFPLA_NET_0_73482, Y => 
        HIEFFPLA_NET_0_73485);
    
    HIEFFPLA_INST_0_57568 : AOI1
      port map(A => \Science_0_exp_packet_0[48]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74808, Y => HIEFFPLA_NET_0_75006);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRY[7]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75301, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[7]\\\\\);
    
    HIEFFPLA_INST_0_70436 : XOR2
      port map(A => HIEFFPLA_NET_0_72159, B => 
        \Timekeeper_0_microseconds[7]\, Y => HIEFFPLA_NET_0_72130);
    
    HIEFFPLA_INST_0_65391 : NOR3B
      port map(A => HIEFFPLA_NET_0_73389, B => 
        HIEFFPLA_NET_0_73276, C => 
        \Science_0/ADC_READ_0/cnt1up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73391);
    
    \Science_0/ADC_READ_0/data_a[5]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[4]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[5]_net_1\);
    
    HIEFFPLA_INST_0_58203 : AND2
      port map(A => \Science_0_exp_packet_0[63]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        Y => HIEFFPLA_NET_0_74830);
    
    HIEFFPLA_INST_0_56360 : XOR2
      port map(A => HIEFFPLA_NET_0_75304, B => 
        HIEFFPLA_NET_0_75295, Y => HIEFFPLA_NET_0_75301);
    
    HIEFFPLA_INST_0_64944 : NOR3A
      port map(A => UC_I2C4_SDA_in, B => 
        \I2C_PassThrough_0.state[3]\, C => 
        \I2C_PassThrough_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73508);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72857, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\);
    
    \Timing_0/s_time[6]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72045, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_time[6]_net_1\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/sda_1\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_72661, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72624, Q => 
        \Sensors_0.Gyro_0.I2C_Master_0.sda_1\);
    
    HIEFFPLA_INST_0_70480 : AND3
      port map(A => \Timekeeper_0_milliseconds[3]\, B => 
        HIEFFPLA_NET_0_72125, C => \Timekeeper_0_milliseconds[4]\, 
        Y => HIEFFPLA_NET_0_72117);
    
    HIEFFPLA_INST_0_65165 : AOI1D
      port map(A => HIEFFPLA_NET_0_73464, B => 
        HIEFFPLA_NET_0_73467, C => HIEFFPLA_NET_0_73428, Y => 
        HIEFFPLA_NET_0_73454);
    
    HIEFFPLA_INST_0_65427 : NAND2
      port map(A => \Science_0/ADC_READ_0/cnt2dn[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2dn[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73380);
    
    HIEFFPLA_INST_0_67300 : AO1
      port map(A => HIEFFPLA_NET_0_72003, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => HIEFFPLA_NET_0_72739, Y => HIEFFPLA_NET_0_72913);
    
    HIEFFPLA_INST_0_66535 : AOI1D
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        C => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73099);
    
    HIEFFPLA_INST_0_59683 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[49]\, B => 
        \Data_Hub_Packets_0_status_packet[53]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74523);
    
    \General_Controller_0/uc_send[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73762, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73601, Q => 
        \General_Controller_0_uc_send[7]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/data_out_1[7]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_72567, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72547, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[7]\);
    
    \Timing_0/s_count[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72023, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_count[2]_net_1\);
    
    HIEFFPLA_INST_0_58996 : NOR3B
      port map(A => HIEFFPLA_NET_0_74469, B => 
        HIEFFPLA_NET_0_74641, C => HIEFFPLA_NET_0_74371, Y => 
        HIEFFPLA_NET_0_74642);
    
    \General_Controller_0/sweep_table_nof_steps[4]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73980, Q => 
        \General_Controller_0/sweep_table_nof_steps[4]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/old_gyro_new_data\ : DFN0P1
      port map(D => \AFLSDF_INV_16\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => 
        \Data_Saving_0/Packet_Saver_0/old_gyro_new_data_i_0\);
    
    HIEFFPLA_INST_0_68464 : AND3C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[3]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[2]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_72645);
    
    HIEFFPLA_INST_0_59585 : MX2
      port map(A => HIEFFPLA_NET_0_74383, B => 
        HIEFFPLA_NET_0_74452, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74534);
    
    \General_Controller_0/sweep_table_step_id[1]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73926, Q => 
        \General_Controller_0/sweep_table_step_id[1]_net_1\);
    
    HIEFFPLA_INST_0_68895 : NOR3B
      port map(A => General_Controller_0_en_sensors, B => 
        HIEFFPLA_NET_0_72528, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, Y
         => HIEFFPLA_NET_0_72529);
    
    HIEFFPLA_INST_0_65353 : XA1B
      port map(A => HIEFFPLA_NET_0_73398, B => 
        \Science_0/ADC_READ_0/cnt1dn[6]_net_1\, C => 
        HIEFFPLA_NET_0_73244, Y => HIEFFPLA_NET_0_73402);
    
    \General_Controller_0/uc_rx_prev_state[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74055, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_prev_state[3]_net_1\);
    
    HIEFFPLA_INST_0_68515 : NAND3
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_i2c_repeat_start\, 
        C => \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72631);
    
    HIEFFPLA_INST_0_57253 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[60]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_75110);
    
    HIEFFPLA_INST_0_70394 : AX1
      port map(A => \Timekeeper_0/old_1MHz_net_1\, B => 
        \s_clks_net_0[4]\, C => \Timekeeper_0_microseconds[0]\, Y
         => HIEFFPLA_NET_0_72151);
    
    HIEFFPLA_INST_0_67832 : AO1A
      port map(A => HIEFFPLA_NET_0_72911, B => 
        HIEFFPLA_NET_0_72749, C => HIEFFPLA_NET_0_72797, Y => 
        HIEFFPLA_NET_0_72791);
    
    HIEFFPLA_INST_0_61396 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[42]\, B => 
        \Timekeeper_0_milliseconds[2]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74204);
    
    HIEFFPLA_INST_0_69762 : AO1A
      port map(A => HIEFFPLA_NET_0_72230, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/isSetup_net_1\, 
        Y => HIEFFPLA_NET_0_72313);
    
    HIEFFPLA_INST_0_65302 : AND3C
      port map(A => HIEFFPLA_NET_0_73416, B => 
        \Science_0/ADC_READ_0/cnt1dn[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt1dn[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73417);
    
    HIEFFPLA_INST_0_58840 : AO1
      port map(A => HIEFFPLA_NET_0_74620, B => 
        HIEFFPLA_NET_0_74372, C => HIEFFPLA_NET_0_74675, Y => 
        HIEFFPLA_NET_0_74676);
    
    HIEFFPLA_INST_0_58092 : AOI1D
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => \Sensors_0_acc_temp[2]\, Y => HIEFFPLA_NET_0_74856);
    
    \General_Controller_0/uc_tx_state[15]\ : DFN1E0P1
      port map(D => HIEFFPLA_NET_0_73573, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[15]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_0[5]\ : DFN0E0C1
      port map(D => 
        \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\);
    
    \Pressure_Signal_Debounce_0/state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73476, CLK => \m_time[7]\, CLR
         => CLKINT_1_Y, Q => 
        \Pressure_Signal_Debounce_0/state[0]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[10]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72803, Q => 
        \Sensors_0_mag_x[10]\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRYSYNC[5]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_11_Q\, 
        CLK => CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[5]\\\\\);
    
    HIEFFPLA_INST_0_57465 : AO1B
      port map(A => \Sensors_0_mag_z[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75037, Y => HIEFFPLA_NET_0_75038);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_new_data\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72287, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        Q => Sensors_0_pressure_new_data);
    
    HIEFFPLA_INST_0_69611 : NOR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        B => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72349);
    
    HIEFFPLA_INST_0_60925 : AND3C
      port map(A => \General_Controller_0/un10_uc_tx_rdy_i[6]\, B
         => \General_Controller_0/un10_uc_tx_rdy_i[7]\, C => 
        \General_Controller_0/un10_uc_tx_rdy_i[5]\, Y => 
        HIEFFPLA_NET_0_74318);
    
    HIEFFPLA_INST_0_58644 : AO1A
      port map(A => HIEFFPLA_NET_0_74655, B => 
        \GS_Readout_0/state[0]_net_1\, C => HIEFFPLA_NET_0_74703, 
        Y => HIEFFPLA_NET_0_74714);
    
    \Timing_0/s_count[7]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72050, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_count[7]_net_1\);
    
    \Science_0/ADC_READ_0/data_b[16]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[16]_net_1\);
    
    HIEFFPLA_INST_0_65199 : AX1C
      port map(A => HIEFFPLA_NET_0_73445, B => 
        \Pressure_Signal_Debounce_0/ms_cnt[6]_net_1\, C => 
        \Pressure_Signal_Debounce_0/ms_cnt[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73447);
    
    HIEFFPLA_INST_0_60360 : MX2
      port map(A => HIEFFPLA_NET_0_74466, B => 
        HIEFFPLA_NET_0_74504, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74427);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[13]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72490, Q => 
        \ch3_data_net_0[9]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[13]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[13]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[13]\);
    
    HIEFFPLA_INST_0_67084 : AO1A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        C => HIEFFPLA_NET_0_72915, Y => HIEFFPLA_NET_0_72968);
    
    HIEFFPLA_INST_0_70126 : AO1A
      port map(A => HIEFFPLA_NET_0_72206, B => 
        HIEFFPLA_NET_0_72275, C => HIEFFPLA_NET_0_72212, Y => 
        HIEFFPLA_NET_0_72213);
    
    HIEFFPLA_INST_0_68608 : AO1E
      port map(A => HIEFFPLA_NET_0_72581, B => 
        HIEFFPLA_NET_0_72582, C => HIEFFPLA_NET_0_72606, Y => 
        HIEFFPLA_NET_0_72607);
    
    HIEFFPLA_INST_0_61915 : OR3A
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => \General_Controller_0/uc_rx_byte[2]_net_1\, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74100);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_2[5]\ : DFN0E0C1
      port map(D => 
        \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\);
    
    HIEFFPLA_INST_0_71116 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_71980, Y => HIEFFPLA_NET_0_75011);
    
    HIEFFPLA_INST_0_67599 : OA1C
      port map(A => HIEFFPLA_NET_0_72957, B => 
        HIEFFPLA_NET_0_72941, C => HIEFFPLA_NET_0_72943, Y => 
        HIEFFPLA_NET_0_72845);
    
    HIEFFPLA_INST_0_65765 : XA1B
      port map(A => HIEFFPLA_NET_0_73293, B => 
        \Science_0/ADC_READ_0/cnt[5]_net_1\, C => 
        HIEFFPLA_NET_0_73241, Y => HIEFFPLA_NET_0_73285);
    
    HIEFFPLA_INST_0_56100 : AO1D
      port map(A => HIEFFPLA_NET_0_75346, B => 
        HIEFFPLA_NET_0_75345, C => 
        \Data_Saving_0/FPGA_Buffer_0/full\, Y => 
        HIEFFPLA_NET_0_75347);
    
    HIEFFPLA_INST_0_55086 : AO1
      port map(A => HIEFFPLA_NET_0_75589, B => 
        HIEFFPLA_NET_0_75585, C => HIEFFPLA_NET_0_75592, Y => 
        HIEFFPLA_NET_0_75594);
    
    HIEFFPLA_INST_0_65019 : XA1
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[6]_net_1\, 
        B => HIEFFPLA_NET_0_73445, C => HIEFFPLA_NET_0_73477, Y
         => HIEFFPLA_NET_0_73487);
    
    \Science_0/ADC_READ_0/data_a[11]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[11]_net_1\);
    
    HIEFFPLA_INST_0_70941 : OA1C
      port map(A => HIEFFPLA_NET_0_72004, B => 
        HIEFFPLA_NET_0_72944, C => HIEFFPLA_NET_0_72831, Y => 
        HIEFFPLA_NET_0_72857);
    
    HIEFFPLA_INST_0_58892 : AND2
      port map(A => \General_Controller_0_gs_id[2]\, B => 
        HIEFFPLA_NET_0_74484, Y => HIEFFPLA_NET_0_74663);
    
    \Science_0/SET_LP_GAIN_0/LA1\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_73182, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73160, Q => LA1_c);
    
    HIEFFPLA_INST_0_64853 : AND3C
      port map(A => HIEFFPLA_NET_0_73600, B => 
        HIEFFPLA_NET_0_73610, C => HIEFFPLA_NET_0_73614, Y => 
        HIEFFPLA_NET_0_73524);
    
    \Science_0/ADC_READ_0/data_a[17]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[17]_net_1\);
    
    HIEFFPLA_INST_0_60969 : AOI1D
      port map(A => \Timekeeper_0_milliseconds[1]\, B => 
        \Timekeeper_0_milliseconds[0]\, C => HIEFFPLA_NET_0_74306, 
        Y => HIEFFPLA_NET_0_74308);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[18]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[18]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[18]\);
    
    HIEFFPLA_INST_0_65423 : AO1E
      port map(A => HIEFFPLA_NET_0_73383, B => 
        HIEFFPLA_NET_0_73385, C => HIEFFPLA_NET_0_73277, Y => 
        HIEFFPLA_NET_0_73381);
    
    HIEFFPLA_INST_0_56748 : AO1
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[1]_net_1\, B => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_75182, Y => HIEFFPLA_NET_0_75216);
    
    HIEFFPLA_INST_0_55261 : AOI1D
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[23]_net_1\, B => 
        \Communications_0/UART_0/rx_clk_count[24]_net_1\, C => 
        \Communications_0/UART_0/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75550);
    
    \General_Controller_0/sweep_table_samples_per_step[9]\ : 
        DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[9]_net_1\);
    
    HIEFFPLA_INST_0_58366 : AO1
      port map(A => \Sensors_0_mag_y[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75103, Y => HIEFFPLA_NET_0_74790);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/num_bytes_1[0]\ : 
        DFN1E1
      port map(D => \AFLSDF_INV_17\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_72549, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_num_bytes[0]\);
    
    HIEFFPLA_INST_0_56642 : MX2
      port map(A => HIEFFPLA_NET_0_75196, B => 
        HIEFFPLA_NET_0_75063, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75229);
    
    HIEFFPLA_INST_0_55292 : AXO5
      port map(A => HIEFFPLA_NET_0_75543, B => 
        \Communications_0/UART_0/tx_state[1]_net_1\, C => 
        \Communications_0/UART_0/tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75544);
    
    \Science_0/ADC_READ_0/cnt[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73288, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73242, Q => 
        \Science_0/ADC_READ_0/cnt[3]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[9]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72807, Q => 
        \Sensors_0_mag_z[9]\);
    
    HIEFFPLA_INST_0_60910 : NOR3B
      port map(A => HIEFFPLA_NET_0_74028, B => 
        HIEFFPLA_NET_0_74319, C => HIEFFPLA_NET_0_74324, Y => 
        HIEFFPLA_NET_0_74321);
    
    \General_Controller_0/sweep_table_sample_skip[14]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[14]_net_1\);
    
    HIEFFPLA_INST_0_66065 : OR3B
      port map(A => \Science_0/DAC_SET_0/cnt[1]_net_1\, B => 
        HIEFFPLA_NET_0_73220, C => 
        \Science_0/DAC_SET_0/cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73221);
    
    HIEFFPLA_INST_0_61747 : AND3
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[1]_net_1\, B
         => \General_Controller_0/sweep_table_sweep_cnt[0]_net_1\, 
        C => 
        \General_Controller_0/sweep_table_sweep_cnt[2]_net_1\, Y
         => HIEFFPLA_NET_0_74148);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72264, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72537, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_59008 : AO1E
      port map(A => HIEFFPLA_NET_0_74360, B => 
        HIEFFPLA_NET_0_74369, C => \GS_Readout_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_74638);
    
    \Science_0/ADC_READ_0/exp_packet_1[26]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[10]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[26]\);
    
    HIEFFPLA_INST_0_67390 : NOR3A
      port map(A => HIEFFPLA_NET_0_72929, B => 
        HIEFFPLA_NET_0_72736, C => HIEFFPLA_NET_0_72739, Y => 
        HIEFFPLA_NET_0_72893);
    
    HIEFFPLA_INST_0_68665 : OA1C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, B
         => HIEFFPLA_NET_0_72664, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72594);
    
    HIEFFPLA_INST_0_68208 : XAI1
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_72706);
    
    HIEFFPLA_INST_0_61054 : AND3
      port map(A => Eject_Signal_Debounce_0_ffu_ejected_out, B
         => \General_Controller_0/flight_state[2]_net_1\, C => 
        HIEFFPLA_NET_0_74249, Y => HIEFFPLA_NET_0_74286);
    
    HIEFFPLA_INST_0_61146 : NAND3C
      port map(A => 
        \General_Controller_0/state_seconds[10]_net_1\, B => 
        \General_Controller_0/state_seconds[19]_net_1\, C => 
        \General_Controller_0/state_seconds[16]_net_1\, Y => 
        HIEFFPLA_NET_0_74264);
    
    HIEFFPLA_INST_0_66510 : NOR3B
      port map(A => HIEFFPLA_NET_0_73064, B => 
        HIEFFPLA_NET_0_73144, C => HIEFFPLA_NET_0_73080, Y => 
        HIEFFPLA_NET_0_73105);
    
    HIEFFPLA_INST_0_59891 : MX2
      port map(A => \Sensors_0_acc_z[5]\, B => 
        \Sensors_0_acc_z[9]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74491);
    
    \GS_Readout_0/wen\ : DFN1E1C1
      port map(D => Communications_0_ext_tx_rdy, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \GS_Readout_0/state[6]_net_1\, Q => GS_Readout_0_wen);
    
    HIEFFPLA_INST_0_67296 : NOR3B
      port map(A => HIEFFPLA_NET_0_72740, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        C => HIEFFPLA_NET_0_72752, Y => HIEFFPLA_NET_0_72915);
    
    \Timekeeper_0/microseconds[15]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72145, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[15]\);
    
    \General_Controller_0/temp_first_byte[7]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73872, Q => 
        \General_Controller_0/temp_first_byte[7]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[12]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72484, Q => 
        \Sensors_0_gyro_y[12]\);
    
    HIEFFPLA_INST_0_55191 : AND2
      port map(A => \Communications_0/UART_0/rx_count[2]_net_1\, 
        B => \Communications_0/UART_0/rx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75563);
    
    HIEFFPLA_INST_0_62004 : AND3C
      port map(A => \General_Controller_0/uc_rx_byte[6]_net_1\, B
         => \General_Controller_0/uc_rx_byte[5]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[7]_net_1\, Y => 
        HIEFFPLA_NET_0_74076);
    
    HIEFFPLA_INST_0_57641 : AO1B
      port map(A => \Sensors_0_gyro_y[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74983, Y => HIEFFPLA_NET_0_74984);
    
    \Timekeeper_0/microseconds[20]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72139, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[20]\);
    
    \Timing_0/m_time[6]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72063, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_time[6]_net_1\);
    
    HIEFFPLA_INST_0_61350 : AX1
      port map(A => HIEFFPLA_NET_0_74261, B => 
        \General_Controller_0/state_seconds[8]_net_1\, C => 
        \General_Controller_0/state_seconds[9]_net_1\, Y => 
        HIEFFPLA_NET_0_74210);
    
    HIEFFPLA_INST_0_66613 : NAND3C
      port map(A => HIEFFPLA_NET_0_73076, B => 
        HIEFFPLA_NET_0_73078, C => HIEFFPLA_NET_0_73082, Y => 
        HIEFFPLA_NET_0_73083);
    
    HIEFFPLA_INST_0_59907 : MX2
      port map(A => HIEFFPLA_NET_0_74535, B => 
        HIEFFPLA_NET_0_74509, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74489);
    
    HIEFFPLA_INST_0_60454 : MX2
      port map(A => HIEFFPLA_NET_0_74558, B => 
        HIEFFPLA_NET_0_74391, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74412);
    
    \EMU_RX_pad/U0/U1\ : IOIN_IB
      port map(YIN => \EMU_RX_pad/U0/NET1\, Y => EMU_RX_c);
    
    HIEFFPLA_INST_0_62941 : XNOR3
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state[3]_net_1\, C => 
        \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73862);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[18]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72282, Q => 
        \Sensors_0_pressure_temp_raw[18]\);
    
    HIEFFPLA_INST_0_67102 : MX2A
      port map(A => HIEFFPLA_NET_0_72917, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[0]\, 
        S => HIEFFPLA_NET_0_72932, Y => HIEFFPLA_NET_0_72963);
    
    HIEFFPLA_INST_0_57318 : AO1
      port map(A => \Science_0_exp_packet_0[16]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74857, Y => HIEFFPLA_NET_0_75078);
    
    HIEFFPLA_INST_0_69777 : OR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[5]_net_1\, 
        C => HIEFFPLA_NET_0_72303, Y => HIEFFPLA_NET_0_72309);
    
    HIEFFPLA_INST_0_62300 : NOR3B
      port map(A => HIEFFPLA_NET_0_74010, B => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, C => 
        \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74011);
    
    HIEFFPLA_INST_0_56078 : XA1A
      port map(A => HIEFFPLA_NET_0_75330, B => 
        HIEFFPLA_NET_0_75262, C => HIEFFPLA_NET_0_75358, Y => 
        HIEFFPLA_NET_0_75353);
    
    HIEFFPLA_INST_0_60503 : MX2
      port map(A => HIEFFPLA_NET_0_74579, B => 
        HIEFFPLA_NET_0_74373, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74404);
    
    HIEFFPLA_INST_0_55056 : NOR3A
      port map(A => \Communications_0/UART_0/rx_count[1]_net_1\, 
        B => \Communications_0/UART_0/rx_count[2]_net_1\, C => 
        \Communications_0/UART_0/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75601);
    
    HIEFFPLA_INST_0_68681 : AND2
      port map(A => \Sensors_0/Gyro_0/L3GD20H_Interface_0_we\, B
         => \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_72589);
    
    HIEFFPLA_INST_0_64801 : AND2
      port map(A => 
        \General_Controller_0/sweep_table_read_wait[31]_net_1\, B
         => HIEFFPLA_NET_0_73815, Y => HIEFFPLA_NET_0_73539);
    
    HIEFFPLA_INST_0_63596 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[10]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_sample_skip[10]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73743);
    
    \Timing_0/m_count[6]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72073, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_count[6]_net_1\);
    
    \General_Controller_0/exp_adc_reset\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74304, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74303, Q => 
        General_Controller_0_exp_adc_reset);
    
    \General_Controller_0/status_bits_1[47]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74199, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[47]\);
    
    HIEFFPLA_INST_0_65082 : AX1C
      port map(A => HIEFFPLA_NET_0_73497, B => 
        \Pressure_Signal_Debounce_0/state[0]_net_1\, C => 
        \Pressure_Signal_Debounce_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73474);
    
    \Sensors_0/Gyro_0/I2C_Master_0/data_out[1]\ : DFN0E1C1
      port map(D => GYRO_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72682, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[1]\);
    
    HIEFFPLA_INST_0_56470 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[7]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[6]\\\\\, C => 
        HIEFFPLA_NET_0_75321, Y => HIEFFPLA_NET_0_75272);
    
    \FMC_DA_pad[4]/U0/U1\ : IOTRI_OB_EB
      port map(D => \FMC_DA_c[4]\, E => \VCC\, DOUT => 
        \FMC_DA_pad[4]/U0/NET1\, EOUT => \FMC_DA_pad[4]/U0/NET2\);
    
    HIEFFPLA_INST_0_67438 : NOR3B
      port map(A => HIEFFPLA_NET_0_72919, B => 
        \Sensors_0/Accelerometer_0/state[8]\, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72881);
    
    HIEFFPLA_INST_0_57581 : AO1
      port map(A => \Sensors_0_pressure_raw[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_75001, Y => HIEFFPLA_NET_0_75002);
    
    HIEFFPLA_INST_0_69985 : NOR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/isSetup_net_1\, 
        C => HIEFFPLA_NET_0_72245, Y => HIEFFPLA_NET_0_72252);
    
    HIEFFPLA_INST_0_69803 : XA1
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[1]_net_1\, 
        C => HIEFFPLA_NET_0_72236, Y => HIEFFPLA_NET_0_72299);
    
    HIEFFPLA_INST_0_65180 : AX1C
      port map(A => HIEFFPLA_NET_0_73443, B => 
        \Pressure_Signal_Debounce_0/ms_cnt[2]_net_1\, C => 
        \Pressure_Signal_Debounce_0/ms_cnt[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73451);
    
    \CU_SYNC_pad/U0/U0\ : IOPAD_IN
      port map(PAD => CU_SYNC, Y => \CU_SYNC_pad/U0/NET1\);
    
    HIEFFPLA_INST_0_69028 : AOI1D
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, B
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        Y => HIEFFPLA_NET_0_72493);
    
    \General_Controller_0/constant_bias_voltage_1[15]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[15]_net_1\);
    
    HIEFFPLA_INST_0_64307 : MX2
      port map(A => HIEFFPLA_NET_0_73727, B => 
        HIEFFPLA_NET_0_73719, S => HIEFFPLA_NET_0_73619, Y => 
        HIEFFPLA_NET_0_73639);
    
    HIEFFPLA_INST_0_60483 : AND2
      port map(A => Communications_0_ext_tx_rdy, B => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74408);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRYSYNC[10]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_6_Q\, CLK
         => CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[10]\\\\\);
    
    HIEFFPLA_INST_0_65937 : AND3C
      port map(A => \Science_0/ADC_READ_0_G3[0]\, B => 
        \Science_0/ADC_READ_0_G3[1]\, C => HIEFFPLA_NET_0_73253, 
        Y => HIEFFPLA_NET_0_73256);
    
    \Science_0/ADC_READ_0/chan2_data[9]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[9]\);
    
    HIEFFPLA_INST_0_63198 : NAND2B
      port map(A => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73810);
    
    \GS_Readout_0/send[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74717, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74630, Q => 
        \GS_Readout_0_send[0]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[2]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72754, Q => 
        \Sensors_0_acc_z[2]\);
    
    \Data_Saving_0/Packet_Saver_0/status_flag\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_74758, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => 
        General_Controller_0_en_data_saving, Q => 
        \Data_Saving_0/Packet_Saver_0/status_flag_net_1\);
    
    HIEFFPLA_INST_0_70293 : AO1A
      port map(A => HIEFFPLA_NET_0_72285, B => 
        \Sensors_0/Pressure_Sensor_0/state[8]\, C => 
        HIEFFPLA_NET_0_72311, Y => HIEFFPLA_NET_0_72180);
    
    HIEFFPLA_INST_0_68870 : NAND3C
      port map(A => HIEFFPLA_NET_0_72485, B => 
        HIEFFPLA_NET_0_72529, C => HIEFFPLA_NET_0_72521, Y => 
        HIEFFPLA_NET_0_72535);
    
    HIEFFPLA_INST_0_67028 : NOR3A
      port map(A => HIEFFPLA_NET_0_72975, B => 
        HIEFFPLA_NET_0_72890, C => HIEFFPLA_NET_0_72913, Y => 
        HIEFFPLA_NET_0_72982);
    
    HIEFFPLA_INST_0_57591 : AO1
      port map(A => \Sensors_0_pressure_raw[12]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74998, Y => HIEFFPLA_NET_0_74999);
    
    \Science_0/ADC_RESET_0/old_enable\ : DFN1E1C1
      port map(D => General_Controller_0_exp_adc_reset, CLK => 
        \s_time[5]\, CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73234, 
        Q => \Science_0/ADC_RESET_0/old_enable_net_1\);
    
    HIEFFPLA_INST_0_62737 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[3]_net_1\, 
        B => HIEFFPLA_NET_0_73884, C => 
        \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73918);
    
    HIEFFPLA_INST_0_59673 : MX2
      port map(A => HIEFFPLA_NET_0_74403, B => 
        HIEFFPLA_NET_0_74423, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74524);
    
    HIEFFPLA_INST_0_70996 : MX2A
      port map(A => HIEFFPLA_NET_0_71994, B => 
        \Science_0/ADC_READ_0_G1[1]\, S => HIEFFPLA_NET_0_73415, 
        Y => HIEFFPLA_NET_0_73265);
    
    HIEFFPLA_INST_0_57977 : AO1
      port map(A => \Science_0_exp_packet_0[28]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74786, Y => HIEFFPLA_NET_0_74889);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[0]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72279, Q => 
        \Sensors_0_pressure_temp_raw[0]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[39]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[5]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[39]\);
    
    HIEFFPLA_INST_0_70210 : AND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72195);
    
    HIEFFPLA_INST_0_68147 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        Y => HIEFFPLA_NET_0_72723);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[2]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72482, Q => 
        \Sensors_0_gyro_y[2]\);
    
    HIEFFPLA_INST_0_68075 : XNOR2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72738);
    
    HIEFFPLA_INST_0_62175 : NOR3B
      port map(A => HIEFFPLA_NET_0_73788, B => 
        HIEFFPLA_NET_0_73900, C => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74036);
    
    \General_Controller_0/sweep_table_read_value[6]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74158, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[6]_net_1\);
    
    \General_Controller_0/constant_bias_voltage_0[2]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[2]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[2]_net_1\);
    
    \Science_0/ADC_READ_0/cnt2dn[0]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73376, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2dn[0]_net_1\);
    
    HIEFFPLA_INST_0_63644 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[10]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_samples_per_point[10]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73735);
    
    HIEFFPLA_INST_0_57384 : AO1
      port map(A => \Sensors_0_gyro_temp[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75060, Y => HIEFFPLA_NET_0_75061);
    
    HIEFFPLA_INST_0_58145 : AO1
      port map(A => \Sensors_0_mag_time[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75147, Y => HIEFFPLA_NET_0_74840);
    
    \General_Controller_0/sweep_table_probe_id[0]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73924, Q => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\);
    
    HIEFFPLA_INST_0_65516 : AND3C
      port map(A => HIEFFPLA_NET_0_73355, B => 
        \Science_0/ADC_READ_0/cnt3dn[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt3dn[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73356);
    
    AFLSDF_INV_4 : INV
      port map(A => \SweepTable_0/WEBP\, Y => \AFLSDF_INV_4\);
    
    \Science_0/SET_LP_GAIN_0/L4WR\ : DFN0C1
      port map(D => \Science_0/SET_LP_GAIN_0/state_i_0[0]\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => L4WR_c);
    
    HIEFFPLA_INST_0_68998 : NOR3B
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, 
        B => HIEFFPLA_NET_0_72502, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        Y => HIEFFPLA_NET_0_72503);
    
    HIEFFPLA_INST_0_68848 : AO1
      port map(A => HIEFFPLA_NET_0_72487, B => 
        \Sensors_0/Gyro_0/I2C_Master_0_write_done\, C => 
        HIEFFPLA_NET_0_72477, Y => HIEFFPLA_NET_0_72541);
    
    HIEFFPLA_INST_0_68221 : AND2B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_72701);
    
    HIEFFPLA_INST_0_70697 : XOR2
      port map(A => \Timing_0/s_time[2]_net_1\, B => 
        HIEFFPLA_NET_0_72033, Y => HIEFFPLA_NET_0_72040);
    
    HIEFFPLA_INST_0_63899 : AO1
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[11]_net_1\, 
        B => HIEFFPLA_NET_0_73579, C => HIEFFPLA_NET_0_73692, Y
         => HIEFFPLA_NET_0_73693);
    
    HIEFFPLA_INST_0_57625 : AO1B
      port map(A => \Sensors_0_acc_x[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74988, Y => HIEFFPLA_NET_0_74989);
    
    HIEFFPLA_INST_0_67873 : AND3C
      port map(A => HIEFFPLA_NET_0_72757, B => 
        HIEFFPLA_NET_0_72776, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72782);
    
    HIEFFPLA_INST_0_64257 : MX2
      port map(A => HIEFFPLA_NET_0_73740, B => 
        HIEFFPLA_NET_0_73732, S => HIEFFPLA_NET_0_73588, Y => 
        HIEFFPLA_NET_0_73644);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[5]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72503, Q => 
        \Sensors_0_gyro_x[5]\);
    
    HIEFFPLA_INST_0_70055 : AND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        C => HIEFFPLA_NET_0_72229, Y => HIEFFPLA_NET_0_72233);
    
    HIEFFPLA_INST_0_55658 : NAND2
      port map(A => \Communications_0/UART_1/rx_count[1]_net_1\, 
        B => \Communications_0/UART_1/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75451);
    
    \Communications_0/UART_0/rx_byte[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75380, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75611, Q => 
        \Communications_0/UART_0/rx_byte[1]_net_1\);
    
    HIEFFPLA_INST_0_70412 : AX1C
      port map(A => \Timekeeper_0_microseconds[17]\, B => 
        HIEFFPLA_NET_0_72162, C => 
        \Timekeeper_0_microseconds[18]\, Y => 
        HIEFFPLA_NET_0_72142);
    
    \General_Controller_0/sweep_table_sample_skip[6]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[6]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[6]_net_1\);
    
    \Science_0/ADC_READ_0/data_b[7]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[7]_net_1\);
    
    HIEFFPLA_INST_0_66598 : MX2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[2]\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[6]\, 
        S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73086);
    
    HIEFFPLA_INST_0_65150 : AND2
      port map(A => \Sensors_0_pressure_raw[16]\, B => 
        \Sensors_0_pressure_raw[18]\, Y => HIEFFPLA_NET_0_73458);
    
    HIEFFPLA_INST_0_70329 : AND2B
      port map(A => HIEFFPLA_NET_0_72267, B => 
        HIEFFPLA_NET_0_72232, Y => HIEFFPLA_NET_0_72173);
    
    HIEFFPLA_INST_0_70264 : NOR3B
      port map(A => \Sensors_0/Pressure_Sensor_0/state[8]\, B => 
        HIEFFPLA_NET_0_72233, C => HIEFFPLA_NET_0_72285, Y => 
        HIEFFPLA_NET_0_72184);
    
    \General_Controller_0/sweep_table_points[5]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[5]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[5]_net_1\);
    
    \General_Controller_0/uc_tx_nextstate[3]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73624, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73857, Q => 
        \General_Controller_0/uc_tx_nextstate[3]_net_1\);
    
    \Communications_0/UART_0/recv[4]\ : DFN1E1C1
      port map(D => \Communications_0/UART_0/rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75551, Q => 
        \Communications_0/UART_0_recv[4]\);
    
    HIEFFPLA_INST_0_68670 : AOI1D
      port map(A => HIEFFPLA_NET_0_72580, B => 
        HIEFFPLA_NET_0_72578, C => HIEFFPLA_NET_0_72662, Y => 
        HIEFFPLA_NET_0_72593);
    
    HIEFFPLA_INST_0_63224 : NOR3A
      port map(A => HIEFFPLA_NET_0_73918, B => 
        HIEFFPLA_NET_0_73786, C => HIEFFPLA_NET_0_73811, Y => 
        HIEFFPLA_NET_0_73802);
    
    HIEFFPLA_INST_0_69413 : AND3A
      port map(A => HIEFFPLA_NET_0_72427, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        C => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72395);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[17]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[17]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[17]\);
    
    HIEFFPLA_INST_0_63116 : NAND3C
      port map(A => HIEFFPLA_NET_0_73848, B => 
        \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        HIEFFPLA_NET_0_73888, Y => HIEFFPLA_NET_0_73825);
    
    HIEFFPLA_INST_0_65942 : MX2
      port map(A => HIEFFPLA_NET_0_73251, B => 
        \Science_0/ADC_READ_0_G3[1]\, S => HIEFFPLA_NET_0_73350, 
        Y => HIEFFPLA_NET_0_73255);
    
    HIEFFPLA_INST_0_65118 : OR2A
      port map(A => \Sensors_0_pressure_raw[11]\, B => 
        HIEFFPLA_NET_0_73466, Y => HIEFFPLA_NET_0_73467);
    
    HIEFFPLA_INST_0_60519 : MX2
      port map(A => HIEFFPLA_NET_0_74451, B => 
        HIEFFPLA_NET_0_74495, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74402);
    
    HIEFFPLA_INST_0_69782 : NAND3
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[1]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72307);
    
    \Science_0/ADC_READ_0/exp_packet_1[15]\ : DFN1E0
      port map(D => \AFLSDF_INV_18\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[15]\);
    
    \Communications_0/UART_0/rx_clk_count[27]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75572, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75554, Q => 
        \Communications_0/UART_0/rx_clk_count[27]_net_1\);
    
    \Science_0/ADC_READ_0/data_a[6]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[5]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[6]_net_1\);
    
    HIEFFPLA_INST_0_59841 : AND2
      port map(A => HIEFFPLA_NET_0_74474, B => 
        HIEFFPLA_NET_0_74371, Y => HIEFFPLA_NET_0_74499);
    
    \Eject_Signal_Debounce_0/old_1kHz\ : DFN1P1
      port map(D => \AFLSDF_INV_19\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => \Eject_Signal_Debounce_0/old_1kHz_i_0\);
    
    \Communications_0/UART_1/tx_clk_count[4]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75407, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_clk_count_i_0[4]\);
    
    \Science_0/DAC_SET_0/old_set\ : DFN1E1C1
      port map(D => \Science_0/SWEEP_SPIDER2_0_SET\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/DAC_SET_0/state[4]_net_1\, Q => 
        \Science_0/DAC_SET_0/old_set_net_1\);
    
    \General_Controller_0/st_ren1\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74175, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74174, Q => 
        General_Controller_0_st_ren1);
    
    HIEFFPLA_INST_0_61152 : NAND3
      port map(A => \General_Controller_0/state_seconds[0]_net_1\, 
        B => \General_Controller_0/state_seconds[1]_net_1\, C => 
        \General_Controller_0/state_seconds[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74262);
    
    HIEFFPLA_INST_0_55599 : AO1C
      port map(A => HIEFFPLA_NET_0_75466, B => 
        HIEFFPLA_NET_0_75475, C => 
        \Communications_0/UART_1/rx_clk_count[27]_net_1\, Y => 
        HIEFFPLA_NET_0_75469);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[4]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72276, Q => \Sensors_0_pressure_raw[4]\);
    
    HIEFFPLA_INST_0_60703 : OR3A
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[2]_net_1\, C => 
        \GS_Readout_0/subState[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74374);
    
    HIEFFPLA_INST_0_55509 : AND3B
      port map(A => HIEFFPLA_NET_0_75451, B => 
        \Communications_0/UART_1/rx_count[2]_net_1\, C => 
        HIEFFPLA_NET_0_75488, Y => HIEFFPLA_NET_0_75493);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[9]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_75244, CLK => CLKINT_0_Y_0, E
         => CLKINT_1_Y, Q => 
        \Data_Saving_0/Interrupt_Generator_0/counter[9]_net_1\);
    
    HIEFFPLA_INST_0_70752 : AND2
      port map(A => HIEFFPLA_NET_0_72019, B => 
        \Timing_0/s_count[6]_net_1\, Y => HIEFFPLA_NET_0_72022);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[5]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72808, Q => 
        \Sensors_0_mag_z[5]\);
    
    \Science_0/DAC_SET_0/vector[11]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73202, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[11]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[24]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[8]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[24]\);
    
    HIEFFPLA_INST_0_55775 : MX2
      port map(A => HIEFFPLA_NET_0_75426, B => 
        HIEFFPLA_NET_0_75425, S => 
        \Communications_0/UART_1/tx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75427);
    
    HIEFFPLA_INST_0_64846 : NOR3A
      port map(A => HIEFFPLA_NET_0_73528, B => 
        HIEFFPLA_NET_0_73522, C => HIEFFPLA_NET_0_73525, Y => 
        HIEFFPLA_NET_0_73526);
    
    HIEFFPLA_INST_0_62775 : OR2A
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73909);
    
    \General_Controller_0/sweep_table_read_value[1]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74163, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[1]_net_1\);
    
    HIEFFPLA_INST_0_64762 : OA1A
      port map(A => \General_Controller_0/uc_tx_state[14]_net_1\, 
        B => HIEFFPLA_NET_0_73558, C => 
        Communications_0_uc_tx_rdy, Y => HIEFFPLA_NET_0_73547);
    
    HIEFFPLA_INST_0_56217 : AX1
      port map(A => \Data_Saving_0/FPGA_Buffer_0/full\, B => 
        \Data_Saving_0/Packet_Saver_0_we\, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[0]\\\\\, Y
         => HIEFFPLA_NET_0_75331);
    
    HIEFFPLA_INST_0_71216 : AXOI2
      port map(A => General_Controller_0_ext_oen, B => 
        \Communications_0/FFU_Command_Checker_0/state[0]_net_1\, 
        C => 
        \Communications_0/FFU_Command_Checker_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_71971);
    
    \General_Controller_0/uc_rx_byte[0]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[0]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte[0]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[3]\ : DFN1E0
      port map(D => \AFLSDF_INV_20\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[3]\);
    
    HIEFFPLA_INST_0_62258 : AND2B
      port map(A => HIEFFPLA_NET_0_73983, B => 
        HIEFFPLA_NET_0_73994, Y => HIEFFPLA_NET_0_74019);
    
    HIEFFPLA_INST_0_59093 : AO1A
      port map(A => HIEFFPLA_NET_0_74597, B => 
        \GS_Readout_0/prevState[0]_net_1\, C => 
        HIEFFPLA_NET_0_74613, Y => HIEFFPLA_NET_0_74614);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73140, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\);
    
    HIEFFPLA_INST_0_68958 : AO1A
      port map(A => HIEFFPLA_NET_0_72475, B => 
        HIEFFPLA_NET_0_72511, C => HIEFFPLA_NET_0_72510, Y => 
        HIEFFPLA_NET_0_72513);
    
    \General_Controller_0/sweep_table_samples_per_point[11]\ : 
        DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[11]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_0[10]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74767, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\);
    
    HIEFFPLA_INST_0_56108 : NOR3B
      port map(A => HIEFFPLA_NET_0_75364, B => 
        HIEFFPLA_NET_0_89700, C => HIEFFPLA_NET_0_75344, Y => 
        HIEFFPLA_NET_0_75345);
    
    HIEFFPLA_INST_0_59133 : NAND3C
      port map(A => HIEFFPLA_NET_0_74585, B => 
        HIEFFPLA_NET_0_74602, C => HIEFFPLA_NET_0_74603, Y => 
        HIEFFPLA_NET_0_74604);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[4]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72783, Q => 
        \Sensors_0_mag_y[4]\);
    
    HIEFFPLA_INST_0_62456 : AND3
      port map(A => HIEFFPLA_NET_0_73775, B => 
        HIEFFPLA_NET_0_74037, C => HIEFFPLA_NET_0_73888, Y => 
        HIEFFPLA_NET_0_73978);
    
    HIEFFPLA_INST_0_61420 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[45]\, B => 
        \Timekeeper_0_milliseconds[5]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74201);
    
    HIEFFPLA_INST_0_65890 : NAND3A
      port map(A => HIEFFPLA_NET_0_73415, B => 
        \Science_0/ADC_READ_0/cnt1up[4]_net_1\, C => 
        HIEFFPLA_NET_0_73276, Y => HIEFFPLA_NET_0_73263);
    
    HIEFFPLA_INST_0_60889 : OR2A
      port map(A => \General_Controller_0/command[6]_net_1\, B
         => \General_Controller_0/command[5]_net_1\, Y => 
        HIEFFPLA_NET_0_74329);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[10]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72800, Q => 
        \Sensors_0_acc_x[10]\);
    
    HIEFFPLA_INST_0_66538 : AND2B
      port map(A => HIEFFPLA_NET_0_73132, B => ACCE_SCL_c, Y => 
        HIEFFPLA_NET_0_73097);
    
    HIEFFPLA_INST_0_55283 : AO1
      port map(A => HIEFFPLA_NET_0_75564, B => 
        HIEFFPLA_NET_0_75545, C => HIEFFPLA_NET_0_75553, Y => 
        HIEFFPLA_NET_0_75546);
    
    HIEFFPLA_INST_0_65123 : NAND2
      port map(A => \Sensors_0_pressure_raw[7]\, B => 
        \Sensors_0_pressure_raw[5]\, Y => HIEFFPLA_NET_0_73465);
    
    \General_Controller_0/uc_rx_state[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73853, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_state[2]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[16]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[16]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[16]\);
    
    HIEFFPLA_INST_0_60140 : MX2
      port map(A => \ch3_data_net_0[11]\, B => 
        \Sensors_0_acc_z[3]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74455);
    
    \Science_0/DAC_SET_0/vector[10]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73203, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[10]_net_1\);
    
    HIEFFPLA_INST_0_65005 : AND2
      port map(A => HIEFFPLA_NET_0_73477, B => 
        HIEFFPLA_NET_0_73482, Y => HIEFFPLA_NET_0_73490);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRY[4]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75292, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[4]\\\\\);
    
    \Timekeeper_0/milliseconds[9]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72093, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[9]\);
    
    HIEFFPLA_INST_0_57311 : AND2
      port map(A => \Sensors_0_gyro_time[17]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75080);
    
    HIEFFPLA_INST_0_66116 : AND2
      port map(A => \Science_0/DAC_SET_0/ADR[0]_net_1\, B => 
        HIEFFPLA_NET_0_73226, Y => HIEFFPLA_NET_0_73204);
    
    HIEFFPLA_INST_0_59000 : NAND2B
      port map(A => \GS_Readout_0/state[5]_net_1\, B => 
        \GS_Readout_0/state[7]_net_1\, Y => HIEFFPLA_NET_0_74640);
    
    HIEFFPLA_INST_0_58115 : AO1
      port map(A => \Sensors_0_mag_y[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_74847, Y => HIEFFPLA_NET_0_74848);
    
    HIEFFPLA_INST_0_63193 : AND3
      port map(A => HIEFFPLA_NET_0_73906, B => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, C => 
        HIEFFPLA_NET_0_73863, Y => HIEFFPLA_NET_0_73812);
    
    HIEFFPLA_INST_0_58400 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[55]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_74779);
    
    AFLSDF_INV_24 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_24\);
    
    HIEFFPLA_INST_0_69118 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[2]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[3]_net_1\, 
        C => HIEFFPLA_NET_0_72556, Y => HIEFFPLA_NET_0_72467);
    
    HIEFFPLA_INST_0_70969 : AX1D
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_71999);
    
    HIEFFPLA_INST_0_68818 : NAND3C
      port map(A => HIEFFPLA_NET_0_72480, B => 
        HIEFFPLA_NET_0_72552, C => HIEFFPLA_NET_0_72498, Y => 
        HIEFFPLA_NET_0_72549);
    
    HIEFFPLA_INST_0_68518 : AND3
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, B => 
        GYRO_SDA_in, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, Y => 
        HIEFFPLA_NET_0_72630);
    
    \GS_Readout_0/prevState[2]\ : DFN1E0C1
      port map(D => \GS_Readout_0/state[2]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \GS_Readout_0/state[6]_net_1\, Q => 
        \GS_Readout_0/prevState[2]_net_1\);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/data_out[5]\ : 
        DFN0E1C1
      port map(D => PRESSURE_SDA_in, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72397, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[5]\);
    
    HIEFFPLA_INST_0_57940 : AOI1
      port map(A => \Sensors_0_pressure_time[13]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_74898, Y => HIEFFPLA_NET_0_74899);
    
    HIEFFPLA_INST_0_70017 : NOR3A
      port map(A => HIEFFPLA_NET_0_72274, B => 
        HIEFFPLA_NET_0_72228, C => HIEFFPLA_NET_0_72231, Y => 
        HIEFFPLA_NET_0_72246);
    
    \General_Controller_0/led2\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74272, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => LED2_c);
    
    \Science_0/ADC_READ_0/chan4_data[6]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[6]\);
    
    HIEFFPLA_INST_0_68393 : NAND3B
      port map(A => HIEFFPLA_NET_0_72650, B => 
        HIEFFPLA_NET_0_72649, C => HIEFFPLA_NET_0_72581, Y => 
        HIEFFPLA_NET_0_72659);
    
    HIEFFPLA_INST_0_63336 : AXO2
      port map(A => HIEFFPLA_NET_0_74015, B => 
        HIEFFPLA_NET_0_74013, C => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73774);
    
    HIEFFPLA_INST_0_63608 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[12]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_sample_skip[12]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73741);
    
    \Communications_0/UART_1/rx_count[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75450, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/rx_count[0]_net_1\);
    
    HIEFFPLA_INST_0_67388 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72894);
    
    HIEFFPLA_INST_0_65041 : NAND3A
      port map(A => CLKINT_1_Y, B => HIEFFPLA_NET_0_73497, C => 
        \Pressure_Signal_Debounce_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73482);
    
    \General_Controller_0/sweep_table_points[7]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[7]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[7]_net_1\);
    
    HIEFFPLA_INST_0_67315 : AOI1C
      port map(A => HIEFFPLA_NET_0_72929, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_72744, Y => HIEFFPLA_NET_0_72909);
    
    HIEFFPLA_INST_0_59336 : MX2
      port map(A => HIEFFPLA_NET_0_74344, B => 
        HIEFFPLA_NET_0_74462, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74566);
    
    HIEFFPLA_INST_0_56276 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[8]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[7]\\\\\, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[6]\\\\\, Y => 
        HIEFFPLA_NET_0_75323);
    
    \Data_Saving_0/Packet_Saver_0/word_cnt[1]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_74753, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[1]_net_1\);
    
    HIEFFPLA_INST_0_59966 : OA1A
      port map(A => HIEFFPLA_NET_0_74432, B => 
        HIEFFPLA_NET_0_74725, C => HIEFFPLA_NET_0_74556, Y => 
        HIEFFPLA_NET_0_74481);
    
    HIEFFPLA_INST_0_65409 : NAND3B
      port map(A => \Science_0/ADC_READ_0/cnt2dn[7]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2dn[6]_net_1\, C => 
        HIEFFPLA_NET_0_73384, Y => HIEFFPLA_NET_0_73385);
    
    HIEFFPLA_INST_0_63578 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[15]_net_1\, B
         => \General_Controller_0/sweep_table_points[15]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73746);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[3]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72801, Q => 
        \Sensors_0_acc_x[3]\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/state[3]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72610, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\);
    
    HIEFFPLA_INST_0_57359 : AO1A
      port map(A => HIEFFPLA_NET_0_75117, B => 
        \Sensors_0_acc_temp[6]\, C => HIEFFPLA_NET_0_75066, Y => 
        HIEFFPLA_NET_0_75067);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[2]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72783, Q => 
        \Sensors_0_mag_y[2]\);
    
    HIEFFPLA_INST_0_66277 : AOI1B
      port map(A => HIEFFPLA_NET_0_73179, B => 
        \Science_0/SET_LP_GAIN_0/state[7]_net_1\, C => 
        HIEFFPLA_NET_0_73156, Y => HIEFFPLA_NET_0_73159);
    
    HIEFFPLA_INST_0_57903 : AO1
      port map(A => \Science_0_exp_packet_0[65]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75133, Y => HIEFFPLA_NET_0_74910);
    
    \General_Controller_0/uc_send[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73766, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73601, Q => 
        \General_Controller_0_uc_send[3]\);
    
    HIEFFPLA_INST_0_69975 : AO1
      port map(A => HIEFFPLA_NET_0_72304, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        C => HIEFFPLA_NET_0_72249, Y => HIEFFPLA_NET_0_72255);
    
    \General_Controller_0/st_waddr[3]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[3]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_waddr[3]\);
    
    \General_Controller_0/state_seconds[14]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74235, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[14]_net_1\);
    
    HIEFFPLA_INST_0_58481 : AND2
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[1]_net_1\, B => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74755);
    
    HIEFFPLA_INST_0_69637 : AO1A
      port map(A => HIEFFPLA_NET_0_72327, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        C => HIEFFPLA_NET_0_72323, Y => HIEFFPLA_NET_0_72339);
    
    HIEFFPLA_INST_0_68803 : NAND2B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, B
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        Y => HIEFFPLA_NET_0_72554);
    
    HIEFFPLA_INST_0_57957 : AO1B
      port map(A => \Sensors_0_pressure_time[15]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, C
         => HIEFFPLA_NET_0_74893, Y => HIEFFPLA_NET_0_74894);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/temp[0]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72907, Q => 
        \Sensors_0_acc_temp[0]\);
    
    HIEFFPLA_INST_0_55940 : XOR2
      port map(A => \Communications_0/UART_1/tx_count[0]_net_1\, 
        B => \Communications_0/UART_1/tx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75389);
    
    HIEFFPLA_INST_0_70755 : AND3
      port map(A => HIEFFPLA_NET_0_72020, B => 
        \Timing_0/s_count[1]_net_1\, C => 
        \Timing_0/s_count[2]_net_1\, Y => HIEFFPLA_NET_0_72021);
    
    HIEFFPLA_INST_0_67729 : AOI1D
      port map(A => HIEFFPLA_NET_0_72842, B => 
        HIEFFPLA_NET_0_72841, C => HIEFFPLA_NET_0_72911, Y => 
        HIEFFPLA_NET_0_72814);
    
    HIEFFPLA_INST_0_62291 : NAND3C
      port map(A => HIEFFPLA_NET_0_74017, B => 
        HIEFFPLA_NET_0_74015, C => HIEFFPLA_NET_0_74000, Y => 
        HIEFFPLA_NET_0_74013);
    
    HIEFFPLA_INST_0_62462 : NOR3A
      port map(A => HIEFFPLA_NET_0_73972, B => 
        HIEFFPLA_NET_0_73786, C => HIEFFPLA_NET_0_73811, Y => 
        HIEFFPLA_NET_0_73977);
    
    HIEFFPLA_INST_0_61299 : AND2
      port map(A => \General_Controller_0/state_seconds[3]_net_1\, 
        B => HIEFFPLA_NET_0_74293, Y => HIEFFPLA_NET_0_74224);
    
    HIEFFPLA_INST_0_58632 : AO1A
      port map(A => HIEFFPLA_NET_0_74655, B => 
        HIEFFPLA_NET_0_74706, C => HIEFFPLA_NET_0_74690, Y => 
        HIEFFPLA_NET_0_74716);
    
    \Data_Saving_0/Packet_Saver_0/data_out[24]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75220, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[24]\);
    
    HIEFFPLA_INST_0_66033 : AND3A
      port map(A => HIEFFPLA_NET_0_73230, B => LDCLK_c, C => 
        \Science_0/DAC_SET_0/cnt[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73231);
    
    HIEFFPLA_INST_0_58129 : AO1
      port map(A => \Sensors_0_mag_time[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75151, Y => HIEFFPLA_NET_0_74844);
    
    HIEFFPLA_INST_0_59201 : NOR3B
      port map(A => HIEFFPLA_NET_0_74662, B => 
        HIEFFPLA_NET_0_74588, C => \GS_Readout_0/state[6]_net_1\, 
        Y => HIEFFPLA_NET_0_74589);
    
    HIEFFPLA_INST_0_59062 : NOR3B
      port map(A => HIEFFPLA_NET_0_74482, B => 
        HIEFFPLA_NET_0_74619, C => HIEFFPLA_NET_0_74459, Y => 
        HIEFFPLA_NET_0_74623);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_2\ : DFN0E0P1
      port map(D => HIEFFPLA_NET_0_73069, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73100, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_2_net_1\);
    
    HIEFFPLA_INST_0_66024 : XOR2
      port map(A => \Science_0/ADC_READ_0/cnt_chan[0]_net_1\, B
         => HIEFFPLA_NET_0_73241, Y => HIEFFPLA_NET_0_73235);
    
    HIEFFPLA_INST_0_54938 : AOI1B
      port map(A => HIEFFPLA_NET_0_75635, B => 
        HIEFFPLA_NET_0_75636, C => HIEFFPLA_NET_0_75629, Y => 
        HIEFFPLA_NET_0_75634);
    
    HIEFFPLA_INST_0_57628 : AOI1
      port map(A => \Science_0_exp_packet_0[47]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74796, Y => HIEFFPLA_NET_0_74988);
    
    HIEFFPLA_INST_0_55328 : MX2C
      port map(A => \Communications_0/UART_0/tx_byte[2]_net_1\, B
         => \Communications_0/UART_0/tx_byte[6]_net_1\, S => 
        \Communications_0/UART_0/tx_count[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75539);
    
    HIEFFPLA_INST_0_57999 : AO1
      port map(A => \Sensors_0_acc_x[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74882, Y => HIEFFPLA_NET_0_74883);
    
    \Science_0/ADC_READ_0/data_a[10]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[10]_net_1\);
    
    HIEFFPLA_INST_0_67046 : OR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[2]\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        Y => HIEFFPLA_NET_0_72980);
    
    HIEFFPLA_INST_0_65113 : AND3C
      port map(A => \Sensors_0_pressure_raw[23]\, B => 
        \Sensors_0_pressure_raw[21]\, C => 
        \Sensors_0_pressure_raw[19]\, Y => HIEFFPLA_NET_0_73468);
    
    \Science_0/ADC_READ_0/exp_packet_1[45]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[11]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[45]\);
    
    \Timekeeper_0/microseconds[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72134, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[3]\);
    
    HIEFFPLA_INST_0_67120 : MX2
      port map(A => HIEFFPLA_NET_0_72892, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[2]\, 
        S => HIEFFPLA_NET_0_72932, Y => HIEFFPLA_NET_0_72961);
    
    HIEFFPLA_INST_0_63406 : MX2
      port map(A => HIEFFPLA_NET_0_73758, B => 
        HIEFFPLA_NET_0_73693, S => HIEFFPLA_NET_0_73608, Y => 
        HIEFFPLA_NET_0_73766);
    
    HIEFFPLA_INST_0_64041 : MX2
      port map(A => HIEFFPLA_NET_0_73640, B => 
        HIEFFPLA_NET_0_73632, S => HIEFFPLA_NET_0_73585, Y => 
        HIEFFPLA_NET_0_73677);
    
    HIEFFPLA_INST_0_62812 : NOR2A
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73896);
    
    HIEFFPLA_INST_0_70415 : XOR2
      port map(A => \Timekeeper_0_microseconds[1]\, B => 
        \Timekeeper_0_microseconds[0]\, Y => HIEFFPLA_NET_0_72140);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRY[1]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75310, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[1]\\\\\);
    
    HIEFFPLA_INST_0_63046 : AO1
      port map(A => HIEFFPLA_NET_0_73835, B => 
        \General_Controller_0/uc_rx_byte[1]_net_1\, C => 
        HIEFFPLA_NET_0_73834, Y => HIEFFPLA_NET_0_73841);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/data_out_1[5]\ : 
        DFN1E1
      port map(D => HIEFFPLA_NET_0_73003, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72795, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[5]\);
    
    HIEFFPLA_INST_0_68353 : NAND3A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72674);
    
    HIEFFPLA_INST_0_70325 : AOI1D
      port map(A => HIEFFPLA_NET_0_72189, B => 
        HIEFFPLA_NET_0_72230, C => HIEFFPLA_NET_0_72194, Y => 
        HIEFFPLA_NET_0_72174);
    
    HIEFFPLA_INST_0_67399 : NAND3C
      port map(A => HIEFFPLA_NET_0_72901, B => CLKINT_1_Y, C => 
        HIEFFPLA_NET_0_72734, Y => HIEFFPLA_NET_0_72891);
    
    HIEFFPLA_INST_0_57535 : AO1
      port map(A => \Sensors_0_acc_z[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74836, Y => HIEFFPLA_NET_0_75017);
    
    HIEFFPLA_INST_0_56176 : XA1
      port map(A => HIEFFPLA_NET_0_75321, B => 
        HIEFFPLA_NET_0_75288, C => HIEFFPLA_NET_0_75326, Y => 
        HIEFFPLA_NET_0_75336);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1E1C0_data_out[2]\\\\/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75285, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \FMC_DA_c[2]\);
    
    HIEFFPLA_INST_0_70490 : AX1C
      port map(A => \Timekeeper_0_milliseconds[11]\, B => 
        HIEFFPLA_NET_0_72119, C => 
        \Timekeeper_0_milliseconds[12]\, Y => 
        HIEFFPLA_NET_0_72113);
    
    \Communications_0/UART_1/rx_state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75436, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/rx_state[0]_net_1\);
    
    HIEFFPLA_INST_0_64507 : AOI1D
      port map(A => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, B => 
        HIEFFPLA_NET_0_73552, C => 
        \General_Controller_0/uc_tx_state[12]_net_1\, Y => 
        HIEFFPLA_NET_0_73611);
    
    HIEFFPLA_INST_0_62935 : NOR3A
      port map(A => HIEFFPLA_NET_0_73900, B => 
        HIEFFPLA_NET_0_73811, C => HIEFFPLA_NET_0_73804, Y => 
        HIEFFPLA_NET_0_73863);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRY[6]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75296, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[6]\\\\\);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[0]\ : DFN1
      port map(D => HIEFFPLA_NET_0_75253, CLK => CLKINT_0_Y_0, Q
         => 
        \Data_Saving_0/Interrupt_Generator_0/counter[0]_net_1\);
    
    HIEFFPLA_INST_0_71066 : AND3
      port map(A => HIEFFPLA_NET_0_74724, B => 
        HIEFFPLA_NET_0_74720, C => 
        \GS_Readout_0/prevState[7]_net_1\, Y => 
        HIEFFPLA_NET_0_71983);
    
    HIEFFPLA_INST_0_69462 : NAND3C
      port map(A => HIEFFPLA_NET_0_72355, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72383);
    
    HIEFFPLA_INST_0_66929 : NAND3C
      port map(A => HIEFFPLA_NET_0_72745, B => 
        HIEFFPLA_NET_0_72921, C => HIEFFPLA_NET_0_72997, Y => 
        HIEFFPLA_NET_0_73002);
    
    HIEFFPLA_INST_0_65288 : NAND2B
      port map(A => HIEFFPLA_NET_0_73421, B => CLKINT_1_Y, Y => 
        HIEFFPLA_NET_0_73422);
    
    \GS_Readout_0/prevState[1]\ : DFN1E0C1
      port map(D => \GS_Readout_0/state[1]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \GS_Readout_0/state[6]_net_1\, Q => 
        \GS_Readout_0/prevState[1]_net_1\);
    
    HIEFFPLA_INST_0_63386 : MX2
      port map(A => HIEFFPLA_NET_0_73760, B => 
        HIEFFPLA_NET_0_73696, S => HIEFFPLA_NET_0_73608, Y => 
        HIEFFPLA_NET_0_73768);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[15]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72484, Q => 
        \Sensors_0_gyro_y[15]\);
    
    \Science_0/ADC_READ_0/chan6_data[10]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[10]\);
    
    HIEFFPLA_INST_0_68058 : MX2
      port map(A => HIEFFPLA_NET_0_72756, B => 
        HIEFFPLA_NET_0_72715, S => HIEFFPLA_NET_0_72876, Y => 
        HIEFFPLA_NET_0_72742);
    
    HIEFFPLA_INST_0_70451 : AND3
      port map(A => \Timekeeper_0_milliseconds[1]\, B => 
        \Timekeeper_0_milliseconds[0]\, C => 
        \Timekeeper_0_milliseconds[2]\, Y => HIEFFPLA_NET_0_72125);
    
    HIEFFPLA_INST_0_68279 : AO1A
      port map(A => GYRO_SCL_c, B => HIEFFPLA_NET_0_72620, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_72691);
    
    HIEFFPLA_INST_0_67775 : AND3
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, C
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72805);
    
    HIEFFPLA_INST_0_57176 : AO1
      port map(A => \Sensors_0_pressure_time[20]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75009, Y => HIEFFPLA_NET_0_75139);
    
    \General_Controller_0/sweep_table_points[2]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[2]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[2]_net_1\);
    
    HIEFFPLA_INST_0_66759 : OR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        B => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73042);
    
    \General_Controller_0/state_seconds[13]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74236, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[13]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/data_out_1[7]\ : 
        DFN1E1
      port map(D => HIEFFPLA_NET_0_73001, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72795, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[7]\);
    
    HIEFFPLA_INST_0_63830 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[1]_net_1\, B
         => 
        \General_Controller_0/sweep_table_sample_skip[1]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73704);
    
    HIEFFPLA_INST_0_70761 : AND3
      port map(A => \Timing_0/s_count[4]_net_1\, B => 
        \Timing_0/s_count[5]_net_1\, C => HIEFFPLA_NET_0_72021, Y
         => HIEFFPLA_NET_0_72019);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/data_out[0]\ : 
        DFN0E1C1
      port map(D => PRESSURE_SDA_in, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72402, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[0]\);
    
    HIEFFPLA_INST_0_70594 : AND3
      port map(A => \s_clks_net_0[9]\, B => 
        \Timing_0/m_time[3]_net_1\, C => HIEFFPLA_NET_0_72069, Y
         => HIEFFPLA_NET_0_72070);
    
    HIEFFPLA_INST_0_57271 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[53]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75100);
    
    HIEFFPLA_INST_0_57781 : AO1
      port map(A => \Sensors_0_pressure_raw[20]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, C
         => HIEFFPLA_NET_0_74943, Y => HIEFFPLA_NET_0_74944);
    
    HIEFFPLA_INST_0_70468 : AND3
      port map(A => \Timekeeper_0_milliseconds[5]\, B => 
        HIEFFPLA_NET_0_72117, C => \Timekeeper_0_milliseconds[6]\, 
        Y => HIEFFPLA_NET_0_72120);
    
    HIEFFPLA_INST_0_66052 : OR3B
      port map(A => HIEFFPLA_NET_0_73213, B => 
        \Science_0/DAC_SET_0/cnt[2]_net_1\, C => 
        HIEFFPLA_NET_0_73223, Y => HIEFFPLA_NET_0_73225);
    
    HIEFFPLA_INST_0_69772 : OR3A
      port map(A => HIEFFPLA_NET_0_72310, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[7]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72311);
    
    HIEFFPLA_INST_0_57245 : AND2
      port map(A => \Sensors_0_gyro_y[12]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75116);
    
    HIEFFPLA_INST_0_68866 : NOR3B
      port map(A => HIEFFPLA_NET_0_72475, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, C
         => \Sensors_0/Gyro_0/I2C_Master_0_s_ack_error\, Y => 
        HIEFFPLA_NET_0_72536);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[1]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72503, Q => 
        \Sensors_0_gyro_x[1]\);
    
    \Science_0/ADC_READ_0/data_b[11]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[11]_net_1\);
    
    HIEFFPLA_INST_0_62131 : OR3A
      port map(A => HIEFFPLA_NET_0_73781, B => 
        HIEFFPLA_NET_0_74154, C => HIEFFPLA_NET_0_73778, Y => 
        HIEFFPLA_NET_0_74045);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72533, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\);
    
    \Science_0/ADC_READ_0/data_b[17]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[17]_net_1\);
    
    HIEFFPLA_INST_0_60689 : MX2
      port map(A => HIEFFPLA_NET_0_74567, B => 
        HIEFFPLA_NET_0_74364, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74376);
    
    \Science_0/ADC_READ_0/chan3_data[2]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[2]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[67]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[11]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[67]\);
    
    HIEFFPLA_INST_0_64504 : AND2B
      port map(A => HIEFFPLA_NET_0_74323, B => 
        \General_Controller_0/un10_uc_tx_rdy_i[1]\, Y => 
        HIEFFPLA_NET_0_73612);
    
    HIEFFPLA_INST_0_57722 : AOI1
      port map(A => \Science_0_exp_packet_0[57]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74821, Y => HIEFFPLA_NET_0_74960);
    
    \Communications_0/UART_1/tx_byte[4]\ : DFN1E1
      port map(D => \General_Controller_0_uc_send[4]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_75385, Q => 
        \Communications_0/UART_1/tx_byte[4]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/data_out_1[6]\ : 
        DFN1E0C1
      port map(D => HIEFFPLA_NET_0_72284, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72270, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[6]\);
    
    HIEFFPLA_INST_0_65844 : MX2
      port map(A => HIEFFPLA_NET_0_73269, B => 
        HIEFFPLA_NET_0_73267, S => 
        \Science_0/ADC_READ_0/chan[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73271);
    
    \ClockDivs_0/cnt_800kHz[0]\ : DFN1C1
      port map(D => \AFLSDF_INV_21\, CLK => CLKINT_0_Y_0, CLR => 
        CLKINT_1_Y, Q => \ClockDivs_0/cnt_800kHz[0]_net_1\);
    
    HIEFFPLA_INST_0_57791 : AO1
      port map(A => \Sensors_0_pressure_raw[21]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, C
         => HIEFFPLA_NET_0_74940, Y => HIEFFPLA_NET_0_74941);
    
    HIEFFPLA_INST_0_68790 : AO1A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        B => HIEFFPLA_NET_0_72479, C => HIEFFPLA_NET_0_72560, Y
         => HIEFFPLA_NET_0_72561);
    
    \Communications_0/UART_0/rx_clk_count[29]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75570, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75554, Q => 
        \Communications_0/UART_0/rx_clk_count[29]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[23]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[23]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[23]\);
    
    \AA_pad/U0/U0\ : IOPAD_IN
      port map(PAD => AA, Y => \AA_pad/U0/NET1\);
    
    \Science_0/ADC_READ_0/cnt[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73284, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73242, Q => 
        \Science_0/ADC_READ_0/cnt[6]_net_1\);
    
    HIEFFPLA_INST_0_62572 : AND3A
      port map(A => HIEFFPLA_NET_0_73810, B => 
        \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73954);
    
    HIEFFPLA_INST_0_67281 : AND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[3]_net_1\, 
        B => CLKINT_1_Y, Y => HIEFFPLA_NET_0_72919);
    
    HIEFFPLA_INST_0_58228 : AO1
      port map(A => \Sensors_0_gyro_x[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74823, Y => HIEFFPLA_NET_0_74824);
    
    HIEFFPLA_INST_0_63293 : NAND3C
      port map(A => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[4]_net_1\, C => 
        \General_Controller_0/uc_rx_substate[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73785);
    
    HIEFFPLA_INST_0_58479 : AOI1
      port map(A => General_Controller_0_status_new_data, B => 
        \Data_Saving_0/Packet_Saver_0/old_status_new_data_i_0\, C
         => \Data_Saving_0/Packet_Saver_0/status_flag_net_1\, Y
         => HIEFFPLA_NET_0_74756);
    
    HIEFFPLA_INST_0_58162 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[15]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75099, Y => HIEFFPLA_NET_0_74836);
    
    HIEFFPLA_INST_0_55245 : AOI1D
      port map(A => HIEFFPLA_NET_0_75580, B => 
        HIEFFPLA_NET_0_75582, C => 
        \Communications_0/UART_0/rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75553);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_3\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[4]\\\\\, CLK => 
        CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_3_Q\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[5]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72800, Q => 
        \Sensors_0_acc_x[5]\);
    
    \Science_0/DAC_SET_0/vector[17]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73196, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[17]_net_1\);
    
    HIEFFPLA_INST_0_67068 : AO1A
      port map(A => HIEFFPLA_NET_0_72971, B => 
        HIEFFPLA_NET_0_72888, C => HIEFFPLA_NET_0_72916, Y => 
        HIEFFPLA_NET_0_72972);
    
    HIEFFPLA_INST_0_60497 : NOR2A
      port map(A => HIEFFPLA_NET_0_74564, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74405);
    
    \Science_0/SET_LP_GAIN_0/old_G2[1]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73172, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/old_G2[1]_net_1\);
    
    HIEFFPLA_INST_0_57988 : NAND2B
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_74886);
    
    HIEFFPLA_INST_0_68405 : MX2
      port map(A => HIEFFPLA_NET_0_72655, B => 
        HIEFFPLA_NET_0_72654, S => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_72657);
    
    HIEFFPLA_INST_0_71164 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[5]\\\\\, B => 
        HIEFFPLA_NET_0_75323, C => HIEFFPLA_NET_0_75260, Y => 
        HIEFFPLA_NET_0_71975);
    
    HIEFFPLA_INST_0_68927 : NAND2A
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0_s_ack_error\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, Y
         => HIEFFPLA_NET_0_72519);
    
    HIEFFPLA_INST_0_60876 : NOR2A
      port map(A => HIEFFPLA_NET_0_74332, B => 
        \General_Controller_0/command[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74333);
    
    HIEFFPLA_INST_0_67291 : AOI1D
      port map(A => HIEFFPLA_NET_0_72898, B => 
        HIEFFPLA_NET_0_72897, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, Y
         => HIEFFPLA_NET_0_72916);
    
    HIEFFPLA_INST_0_62729 : AOI1B
      port map(A => HIEFFPLA_NET_0_73937, B => 
        HIEFFPLA_NET_0_73919, C => HIEFFPLA_NET_0_74035, Y => 
        HIEFFPLA_NET_0_73920);
    
    HIEFFPLA_INST_0_61107 : AND2B
      port map(A => \Timekeeper_0_milliseconds[14]\, B => 
        \Timekeeper_0_milliseconds[10]\, Y => 
        HIEFFPLA_NET_0_74275);
    
    HIEFFPLA_INST_0_66806 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        B => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73031);
    
    \Science_0/DAC_SET_0/cnt[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73215, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/cnt[4]_net_1\);
    
    HIEFFPLA_INST_0_68963 : AOI1D
      port map(A => General_Controller_0_en_sensors, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, C
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72512);
    
    HIEFFPLA_INST_0_57209 : AO1
      port map(A => \Sensors_0_pressure_time[12]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75089, Y => HIEFFPLA_NET_0_75129);
    
    HIEFFPLA_INST_0_68731 : XOR2
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, B => 
        HIEFFPLA_NET_0_72634, Y => HIEFFPLA_NET_0_72575);
    
    \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_1\ : DFN0E0P1
      port map(D => HIEFFPLA_NET_0_72643, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72619, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_1_net_1\);
    
    HIEFFPLA_INST_0_57223 : AND2
      port map(A => \Sensors_0_pressure_raw[23]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, Y
         => HIEFFPLA_NET_0_75122);
    
    HIEFFPLA_INST_0_66604 : MX2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[0]\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[5]\, 
        S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73085);
    
    HIEFFPLA_INST_0_62022 : XA1B
      port map(A => 
        \General_Controller_0/uc_rx_prev_state[4]_net_1\, B => 
        \General_Controller_0/uc_rx_prev_state[3]_net_1\, C => 
        Communications_0_uc_rx_rdy, Y => HIEFFPLA_NET_0_74069);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[11]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72803, Q => 
        \Sensors_0_mag_x[11]\);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_16\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[6]\\\\\, CLK => 
        CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_16_Q\);
    
    HIEFFPLA_INST_0_65299 : NOR3A
      port map(A => \Science_0/ADC_READ_0/newflag_net_1\, B => 
        \Science_0/ADC_READ_0/chan[0]_net_1\, C => 
        \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73418);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/isSetup\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72559, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/isSetup_net_1\);
    
    HIEFFPLA_INST_0_59869 : MX2
      port map(A => \Science_0_chan3_data[0]\, B => 
        \Science_0_chan3_data[4]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74494);
    
    HIEFFPLA_INST_0_56485 : AX1
      port map(A => \Data_Saving_0/FPGA_Buffer_0/empty\, B => 
        FMC_NOE_c, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[0]\\\\\, Y
         => HIEFFPLA_NET_0_75268);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_1\ : 
        DFN0E0P1
      port map(D => HIEFFPLA_NET_0_72362, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72384, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_1_net_1\);
    
    HIEFFPLA_INST_0_70342 : AOI1D
      port map(A => General_Controller_0_st_ren1, B => 
        \SweepTable_0/WEBP\, C => 
        \General_Controller_0_st_raddr_1[3]\, Y => 
        \TableSelect_0_RADDR[3]\);
    
    HIEFFPLA_INST_0_62120 : NOR2A
      port map(A => HIEFFPLA_NET_0_73943, B => 
        \General_Controller_0/uc_rx_prev_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74048);
    
    \ACCE_SCL_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => ACCE_SCL_c, E => \VCC\, DOUT => 
        \ACCE_SCL_pad/U0/NET1\, EOUT => \ACCE_SCL_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_66122 : MX2B
      port map(A => \Science_0/DAC_SET_0/vector[10]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73202);
    
    HIEFFPLA_INST_0_63967 : MX2
      port map(A => HIEFFPLA_NET_0_73655, B => 
        HIEFFPLA_NET_0_73647, S => HIEFFPLA_NET_0_73599, Y => 
        HIEFFPLA_NET_0_73684);
    
    HIEFFPLA_INST_0_62613 : AO1
      port map(A => HIEFFPLA_NET_0_73917, B => 
        HIEFFPLA_NET_0_73775, C => HIEFFPLA_NET_0_73878, Y => 
        HIEFFPLA_NET_0_73945);
    
    HIEFFPLA_INST_0_61808 : NOR3B
      port map(A => HIEFFPLA_NET_0_74124, B => 
        HIEFFPLA_NET_0_73780, C => HIEFFPLA_NET_0_73786, Y => 
        HIEFFPLA_NET_0_74125);
    
    HIEFFPLA_INST_0_61508 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[56]\, B => 
        \Timekeeper_0_milliseconds[16]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74190);
    
    HIEFFPLA_INST_0_61412 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[44]\, B => 
        \Timekeeper_0_milliseconds[4]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74202);
    
    \Data_Saving_0/Packet_Saver_0/data_out[18]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75227, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[18]\);
    
    HIEFFPLA_INST_0_62853 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state[1]_net_1\, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73881);
    
    HIEFFPLA_INST_0_59256 : MX2
      port map(A => \Science_0_chan4_data[6]\, B => 
        \Science_0_chan4_data[10]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74579);
    
    HIEFFPLA_INST_0_58346 : AO1
      port map(A => \Sensors_0_gyro_x[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74795, Y => HIEFFPLA_NET_0_74796);
    
    \Communications_0/UART_1/tx_state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75384, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_state[0]_net_1\);
    
    HIEFFPLA_INST_0_56493 : AX1C
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[1]\\\\\, B
         => HIEFFPLA_NET_0_75369, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[2]\\\\\, Y
         => HIEFFPLA_NET_0_75265);
    
    HIEFFPLA_INST_0_69400 : NOR3B
      port map(A => HIEFFPLA_NET_0_72351, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        C => HIEFFPLA_NET_0_72394, Y => HIEFFPLA_NET_0_72398);
    
    HIEFFPLA_INST_0_68327 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, B => 
        HIEFFPLA_NET_0_72678, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72681);
    
    HIEFFPLA_INST_0_69455 : MX2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_72383, S => PRESSURE_SCL_c, Y => 
        HIEFFPLA_NET_0_72384);
    
    HIEFFPLA_INST_0_64227 : MX2
      port map(A => HIEFFPLA_NET_0_73743, B => 
        HIEFFPLA_NET_0_73735, S => HIEFFPLA_NET_0_73588, Y => 
        HIEFFPLA_NET_0_73647);
    
    HIEFFPLA_INST_0_60318 : MX2
      port map(A => HIEFFPLA_NET_0_74392, B => 
        HIEFFPLA_NET_0_74576, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74432);
    
    HIEFFPLA_INST_0_68183 : AX1C
      port map(A => HIEFFPLA_NET_0_72711, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72712);
    
    HIEFFPLA_INST_0_69257 : AND3B
      port map(A => HIEFFPLA_NET_0_72436, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, Y
         => HIEFFPLA_NET_0_72437);
    
    HIEFFPLA_INST_0_66111 : OA1A
      port map(A => \Science_0/SWEEP_SPIDER2_0_SET\, B => 
        \Science_0/DAC_SET_0/old_set_net_1\, C => 
        \Science_0/DAC_SET_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73207);
    
    HIEFFPLA_INST_0_64810 : AX1C
      port map(A => HIEFFPLA_NET_0_73780, B => 
        HIEFFPLA_NET_0_74013, C => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73536);
    
    HIEFFPLA_INST_0_61789 : AX1C
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[5]_net_1\, B
         => HIEFFPLA_NET_0_74150, C => 
        \General_Controller_0/sweep_table_sweep_cnt[6]_net_1\, Y
         => HIEFFPLA_NET_0_74132);
    
    HIEFFPLA_INST_0_55322 : MX2C
      port map(A => \Communications_0/UART_0/tx_byte[0]_net_1\, B
         => \Communications_0/UART_0/tx_byte[4]_net_1\, S => 
        \Communications_0/UART_0/tx_count[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75540);
    
    \FMC_DA_pad[0]/U0/U1\ : IOTRI_OB_EB
      port map(D => \FMC_DA_c[0]\, E => \VCC\, DOUT => 
        \FMC_DA_pad[0]/U0/NET1\, EOUT => \FMC_DA_pad[0]/U0/NET2\);
    
    HIEFFPLA_INST_0_70387 : AND2
      port map(A => HIEFFPLA_NET_0_72160, B => 
        \Timekeeper_0_microseconds[21]\, Y => 
        HIEFFPLA_NET_0_72153);
    
    HIEFFPLA_INST_0_68647 : NOR3A
      port map(A => HIEFFPLA_NET_0_72702, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, C => 
        HIEFFPLA_NET_0_72591, Y => HIEFFPLA_NET_0_72597);
    
    HIEFFPLA_INST_0_58110 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_74851);
    
    \Communications_0/FFU_Command_Checker_0/state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75623, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/FFU_Command_Checker_0/state[0]_net_1\);
    
    HIEFFPLA_INST_0_58106 : AO1
      port map(A => \Science_0_exp_packet_0[15]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_75118, Y => HIEFFPLA_NET_0_74853);
    
    HIEFFPLA_INST_0_88377 : XNOR3
      port map(A => HIEFFPLA_NET_0_88381, B => 
        HIEFFPLA_NET_0_75304, C => HIEFFPLA_NET_0_75320, Y => 
        HIEFFPLA_NET_0_89700);
    
    \Data_Saving_0/Packet_Saver_0/packet_select[10]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74767, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\);
    
    AFLSDF_INV_5 : INV
      port map(A => CLKINT_1_Y, Y => \AFLSDF_INV_5\);
    
    HIEFFPLA_INST_0_56881 : MX2
      port map(A => HIEFFPLA_NET_0_74999, B => 
        HIEFFPLA_NET_0_74927, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75200);
    
    HIEFFPLA_INST_0_58201 : AO1
      port map(A => \Sensors_0_acc_time[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74830, Y => HIEFFPLA_NET_0_74831);
    
    HIEFFPLA_INST_0_60856 : NAND2B
      port map(A => HIEFFPLA_NET_0_74327, B => 
        HIEFFPLA_NET_0_74334, Y => HIEFFPLA_NET_0_74339);
    
    HIEFFPLA_INST_0_55627 : XA1
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[26]_net_1\, B => 
        HIEFFPLA_NET_0_75470, C => HIEFFPLA_NET_0_75437, Y => 
        HIEFFPLA_NET_0_75461);
    
    HIEFFPLA_INST_0_63680 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[0]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_nof_steps[0]_net_1\, S
         => \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73729);
    
    HIEFFPLA_INST_0_70159 : OR3B
      port map(A => HIEFFPLA_NET_0_72242, B => 
        HIEFFPLA_NET_0_72275, C => HIEFFPLA_NET_0_72191, Y => 
        HIEFFPLA_NET_0_72205);
    
    HIEFFPLA_INST_0_68027 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        B => \Sensors_0/Accelerometer_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72749);
    
    \General_Controller_0/gs_id[5]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73922, Q => 
        \General_Controller_0_gs_id[5]\);
    
    HIEFFPLA_INST_0_65538 : AOI1B
      port map(A => HIEFFPLA_NET_0_73356, B => 
        HIEFFPLA_NET_0_73353, C => HIEFFPLA_NET_0_73277, Y => 
        HIEFFPLA_NET_0_73349);
    
    HIEFFPLA_INST_0_58417 : AOI1
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/old_gyro_new_data_i_0\, B
         => Sensors_0_gyro_new_data, C => 
        \Data_Saving_0/Packet_Saver_0/gyro_flag_net_1\, Y => 
        HIEFFPLA_NET_0_74773);
    
    HIEFFPLA_INST_0_66695 : AND3C
      port map(A => HIEFFPLA_NET_0_73058, B => 
        HIEFFPLA_NET_0_73066, C => HIEFFPLA_NET_0_73110, Y => 
        HIEFFPLA_NET_0_73061);
    
    HIEFFPLA_INST_0_61138 : AND2
      port map(A => \s_clks_net_0[18]\, B => 
        \General_Controller_0/old_status_packet_clk_i_0\, Y => 
        HIEFFPLA_NET_0_74267);
    
    HIEFFPLA_INST_0_66903 : AO1A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        C => HIEFFPLA_NET_0_72861, Y => HIEFFPLA_NET_0_73008);
    
    HIEFFPLA_INST_0_66463 : AO1A
      port map(A => ACCE_SCL_c, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        C => HIEFFPLA_NET_0_73051, Y => HIEFFPLA_NET_0_73114);
    
    HIEFFPLA_INST_0_65325 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt1dn[0]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt1dn[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt1dn[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73410);
    
    HIEFFPLA_INST_0_70633 : AND3
      port map(A => HIEFFPLA_NET_0_72059, B => 
        \Timing_0/s_count[1]_net_1\, C => HIEFFPLA_NET_0_72057, Y
         => HIEFFPLA_NET_0_72058);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_WADDR[5]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75291, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\);
    
    \Communications_0/UART_0/tx_byte[1]\ : DFN1E1
      port map(D => \GS_Readout_0_send[1]\, CLK => CLKINT_0_Y_0, 
        E => HIEFFPLA_NET_0_75504, Q => 
        \Communications_0/UART_0/tx_byte[1]_net_1\);
    
    HIEFFPLA_INST_0_63764 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[6]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[6]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73715);
    
    HIEFFPLA_INST_0_60952 : AO1
      port map(A => HIEFFPLA_NET_0_74311, B => 
        \General_Controller_0/flight_state[4]_net_1\, C => 
        HIEFFPLA_NET_0_74309, Y => HIEFFPLA_NET_0_74312);
    
    HIEFFPLA_INST_0_67628 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        B => General_Controller_0_en_sensors, Y => 
        HIEFFPLA_NET_0_72839);
    
    \General_Controller_0/uc_rx_state_0[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73867, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\);
    
    \Timekeeper_0/milliseconds[19]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72106, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[19]\);
    
    HIEFFPLA_INST_0_68477 : AO1A
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, 
        B => HIEFFPLA_NET_0_72620, C => HIEFFPLA_NET_0_72626, Y
         => HIEFFPLA_NET_0_72641);
    
    HIEFFPLA_INST_0_57156 : AND2
      port map(A => \Sensors_0_pressure_time[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, Y
         => HIEFFPLA_NET_0_75149);
    
    CLKINT_0 : CLKINT
      port map(A => CLOCK_c, Y => CLKINT_0_Y_0);
    
    HIEFFPLA_INST_0_57289 : AND2
      port map(A => \Sensors_0_gyro_time[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75091);
    
    HIEFFPLA_INST_0_61721 : AND3
      port map(A => HIEFFPLA_NET_0_73779, B => 
        \General_Controller_0/sweep_table_read_wait[30]_net_1\, C
         => 
        \General_Controller_0/sweep_table_read_wait[31]_net_1\, Y
         => HIEFFPLA_NET_0_74154);
    
    HIEFFPLA_INST_0_66184 : AO1B
      port map(A => \Science_0/SET_LP_GAIN_0/state[6]_net_1\, B
         => \Science_0/ADC_READ_0_G2[0]\, C => 
        HIEFFPLA_NET_0_73184, Y => HIEFFPLA_NET_0_73185);
    
    HIEFFPLA_INST_0_63067 : NAND3C
      port map(A => HIEFFPLA_NET_0_73824, B => 
        HIEFFPLA_NET_0_73822, C => HIEFFPLA_NET_0_73820, Y => 
        HIEFFPLA_NET_0_73836);
    
    HIEFFPLA_INST_0_57066 : MX2
      port map(A => HIEFFPLA_NET_0_74947, B => 
        HIEFFPLA_NET_0_74886, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75173);
    
    HIEFFPLA_INST_0_65601 : NOR3B
      port map(A => HIEFFPLA_NET_0_73331, B => 
        HIEFFPLA_NET_0_73276, C => 
        \Science_0/ADC_READ_0/cnt3up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73333);
    
    HIEFFPLA_INST_0_57251 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[58]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_75112);
    
    HIEFFPLA_INST_0_55579 : NOR2A
      port map(A => \Communications_0/UART_1/rx_state[1]_net_1\, 
        B => \Communications_0/UART_1/rx_clk_count[26]_net_1\, Y
         => HIEFFPLA_NET_0_75476);
    
    HIEFFPLA_INST_0_60971 : AO1A
      port map(A => HIEFFPLA_NET_0_74313, B => 
        HIEFFPLA_NET_0_74305, C => 
        General_Controller_0_en_sensors, Y => 
        HIEFFPLA_NET_0_74307);
    
    \Data_Saving_0/Packet_Saver_0/data_out[13]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75232, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[13]\);
    
    HIEFFPLA_INST_0_56461 : OR2A
      port map(A => HIEFFPLA_NET_0_75276, B => 
        HIEFFPLA_NET_0_75331, Y => HIEFFPLA_NET_0_75275);
    
    HIEFFPLA_INST_0_62341 : NOR3B
      port map(A => HIEFFPLA_NET_0_74083, B => 
        HIEFFPLA_NET_0_73881, C => HIEFFPLA_NET_0_74093, Y => 
        HIEFFPLA_NET_0_74002);
    
    HIEFFPLA_INST_0_68052 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        Y => HIEFFPLA_NET_0_72745);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRYSYNC[8]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_19_Q\, 
        CLK => CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[8]\\\\\);
    
    HIEFFPLA_INST_0_70026 : NAND3C
      port map(A => HIEFFPLA_NET_0_72237, B => 
        HIEFFPLA_NET_0_72223, C => HIEFFPLA_NET_0_72222, Y => 
        HIEFFPLA_NET_0_72243);
    
    \Sensors_0/Gyro_0/I2C_Master_0/state[4]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72609, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\);
    
    \General_Controller_0/sweep_table_samples_per_step[11]\ : 
        DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[11]_net_1\);
    
    HIEFFPLA_INST_0_71016 : AO1A
      port map(A => \General_Controller_0/uc_tx_state[0]_net_1\, 
        B => HIEFFPLA_NET_0_71987, C => HIEFFPLA_NET_0_73552, Y
         => HIEFFPLA_NET_0_73528);
    
    HIEFFPLA_INST_0_68150 : NAND3C
      port map(A => HIEFFPLA_NET_0_72720, B => 
        HIEFFPLA_NET_0_72796, C => HIEFFPLA_NET_0_72781, Y => 
        HIEFFPLA_NET_0_72721);
    
    HIEFFPLA_INST_0_70578 : XA1B
      port map(A => HIEFFPLA_NET_0_72031, B => 
        \Timing_0/m_count[5]_net_1\, C => HIEFFPLA_NET_0_72083, Y
         => HIEFFPLA_NET_0_72074);
    
    HIEFFPLA_INST_0_69616 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72345);
    
    HIEFFPLA_INST_0_66001 : NAND2B
      port map(A => \Science_0/ADC_READ_0/state[1]_net_1\, B => 
        HIEFFPLA_NET_0_73241, Y => HIEFFPLA_NET_0_73242);
    
    \Science_0/ADC_READ_0/cnt3dn[2]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73345, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3dn[2]_net_1\);
    
    HIEFFPLA_INST_0_69213 : NAND3B
      port map(A => HIEFFPLA_NET_0_72554, B => 
        HIEFFPLA_NET_0_72435, C => HIEFFPLA_NET_0_72488, Y => 
        HIEFFPLA_NET_0_72445);
    
    HIEFFPLA_INST_0_58413 : OA1C
      port map(A => HIEFFPLA_NET_0_74775, B => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, C => 
        HIEFFPLA_NET_0_74773, Y => HIEFFPLA_NET_0_74774);
    
    \Science_0/ADC_READ_0/chan4_data[11]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[17]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[11]\);
    
    HIEFFPLA_INST_0_57299 : AND2
      port map(A => \Sensors_0_pressure_raw[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75085);
    
    HIEFFPLA_INST_0_67282 : NOR2A
      port map(A => HIEFFPLA_NET_0_72935, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, Y
         => HIEFFPLA_NET_0_72918);
    
    HIEFFPLA_INST_0_65870 : MX2
      port map(A => \Science_0/ADC_READ_0_G2[1]\, B => 
        \Science_0/ADC_READ_0_G4[1]\, S => 
        \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73267);
    
    \Communications_0/UART_1/tx_byte[6]\ : DFN1E1
      port map(D => \General_Controller_0_uc_send[6]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_75385, Q => 
        \Communications_0/UART_1/tx_byte[6]_net_1\);
    
    HIEFFPLA_INST_0_70007 : NOR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_s_ack_error\, B
         => HIEFFPLA_NET_0_72275, C => HIEFFPLA_NET_0_72246, Y
         => HIEFFPLA_NET_0_72248);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/data_out[5]\ : 
        DFN0E1C1
      port map(D => ACCE_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73119, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\);
    
    HIEFFPLA_INST_0_66637 : NAND2A
      port map(A => HIEFFPLA_NET_0_73132, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_repeat_start\, 
        Y => HIEFFPLA_NET_0_73077);
    
    HIEFFPLA_INST_0_68733 : NOR2A
      port map(A => HIEFFPLA_NET_0_72634, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_72574);
    
    \Communications_0/UART_1/recv[4]\ : DFN1E1C1
      port map(D => \Communications_0/UART_1/rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75441, Q => \Communications_0_uc_recv[4]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[16]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[0]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[16]\);
    
    \UC_UART_RX_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => UC_UART_RX_c, E => \VCC\, DOUT => 
        \UC_UART_RX_pad/U0/NET1\, EOUT => 
        \UC_UART_RX_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_67228 : AND2
      port map(A => HIEFFPLA_NET_0_72872, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72934);
    
    HIEFFPLA_INST_0_55547 : MX2A
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\, B => 
        HIEFFPLA_NET_0_75469, S => HIEFFPLA_NET_0_75480, Y => 
        HIEFFPLA_NET_0_75482);
    
    \Communications_0/UART_1/rx_byte[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75378, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75492, Q => 
        \Communications_0/UART_1/rx_byte[4]_net_1\);
    
    \Timing_0/s_count[6]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72051, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_count[6]_net_1\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/data_out_rdy\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_73051, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73114, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\);
    
    HIEFFPLA_INST_0_69343 : OA1A
      port map(A => HIEFFPLA_NET_0_72412, B => PRESSURE_SCL_c, C
         => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72414);
    
    \Timing_0/m_count[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72079, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_count[2]_net_1\);
    
    HIEFFPLA_INST_0_68066 : AO1C
      port map(A => HIEFFPLA_NET_0_72734, B => 
        HIEFFPLA_NET_0_72744, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, Y
         => HIEFFPLA_NET_0_72741);
    
    HIEFFPLA_INST_0_55017 : XO1
      port map(A => \General_Controller_0_unit_id[3]\, B => 
        \Communications_0/UART_0_recv[3]\, C => 
        HIEFFPLA_NET_0_75621, Y => HIEFFPLA_NET_0_75615);
    
    HIEFFPLA_INST_0_67426 : AO1D
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        C => HIEFFPLA_NET_0_72761, Y => HIEFFPLA_NET_0_72884);
    
    \General_Controller_0/sweep_table_sample_skip[12]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[12]_net_1\);
    
    \General_Controller_0/sweep_table_read_value[10]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74169, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[10]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72859, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\);
    
    HIEFFPLA_INST_0_66837 : AOI1A
      port map(A => HIEFFPLA_NET_0_73098, B => 
        HIEFFPLA_NET_0_73108, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73024);
    
    \Science_0/ADC_READ_0/data_b[1]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[0]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[1]_net_1\);
    
    HIEFFPLA_INST_0_63632 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[8]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[8]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73737);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/temp[6]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72555, Q => 
        \Sensors_0_gyro_temp[6]\);
    
    HIEFFPLA_INST_0_66168 : NOR2A
      port map(A => \Science_0/DAC_SET_0/vector[4]_net_1\, B => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73191);
    
    HIEFFPLA_INST_0_59475 : AO1
      port map(A => HIEFFPLA_NET_0_74445, B => 
        HIEFFPLA_NET_0_74341, C => HIEFFPLA_NET_0_74505, Y => 
        HIEFFPLA_NET_0_74549);
    
    \UC_UART_TX_pad/U0/U0\ : IOPAD_IN
      port map(PAD => UC_UART_TX, Y => \UC_UART_TX_pad/U0/NET1\);
    
    \Science_0/ADC_READ_0/chan5_data[6]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[6]\);
    
    HIEFFPLA_INST_0_67510 : NOR3B
      port map(A => HIEFFPLA_NET_0_72740, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        C => HIEFFPLA_NET_0_72752, Y => HIEFFPLA_NET_0_72861);
    
    \Science_0/ADC_READ_0/chan1_data[3]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[3]\);
    
    HIEFFPLA_INST_0_57428 : AO1
      port map(A => \Sensors_0_gyro_temp[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74873, Y => HIEFFPLA_NET_0_75049);
    
    \General_Controller_0/sweep_table_points[3]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[3]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[3]_net_1\);
    
    HIEFFPLA_INST_0_70418 : XOR2
      port map(A => HIEFFPLA_NET_0_72160, B => 
        \Timekeeper_0_microseconds[21]\, Y => 
        HIEFFPLA_NET_0_72138);
    
    HIEFFPLA_INST_0_56929 : MX2
      port map(A => HIEFFPLA_NET_0_74981, B => 
        HIEFFPLA_NET_0_74909, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75194);
    
    \Science_0/ADC_READ_0/cnt1dn[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73405, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1dn[3]_net_1\);
    
    HIEFFPLA_INST_0_60385 : MX2
      port map(A => \Science_0_chan7_data[1]\, B => 
        \Science_0_chan7_data[5]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74423);
    
    HIEFFPLA_INST_0_67769 : NAND3C
      port map(A => HIEFFPLA_NET_0_72930, B => 
        HIEFFPLA_NET_0_72785, C => HIEFFPLA_NET_0_72768, Y => 
        HIEFFPLA_NET_0_72806);
    
    HIEFFPLA_INST_0_58546 : NAND3C
      port map(A => \Eject_Signal_Debounce_0/state[0]_net_1\, B
         => HIEFFPLA_NET_0_74739, C => HIEFFPLA_NET_0_74736, Y
         => HIEFFPLA_NET_0_74738);
    
    HIEFFPLA_INST_0_70573 : AOI1B
      port map(A => HIEFFPLA_NET_0_72082, B => 
        HIEFFPLA_NET_0_72081, C => HIEFFPLA_NET_0_72075, Y => 
        HIEFFPLA_NET_0_72076);
    
    HIEFFPLA_INST_0_64337 : MX2
      port map(A => HIEFFPLA_NET_0_73724, B => 
        HIEFFPLA_NET_0_73716, S => HIEFFPLA_NET_0_73619, Y => 
        HIEFFPLA_NET_0_73636);
    
    HIEFFPLA_INST_0_62149 : NOR3A
      port map(A => HIEFFPLA_NET_0_73897, B => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74042);
    
    \Science_0/ADC_READ_0/exp_packet_1[23]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[7]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[23]\);
    
    \I2C_PassThrough_0/cnt[0]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73505, CLK => CLKINT_0_Y_0, Q
         => \I2C_PassThrough_0/cnt[0]_net_1\);
    
    HIEFFPLA_INST_0_65670 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt4dn[5]_net_1\, B => 
        HIEFFPLA_NET_0_73322, C => HIEFFPLA_NET_0_73274, Y => 
        HIEFFPLA_NET_0_73313);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[9]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72803, Q => 
        \Sensors_0_mag_x[9]\);
    
    HIEFFPLA_INST_0_58466 : OR3A
      port map(A => General_Controller_0_en_data_saving, B => 
        HIEFFPLA_NET_0_74759, C => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74760);
    
    \Science_0/ADC_READ_0/chan4_data[0]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[0]\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_WADDR[8]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75295, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[8]\\\\\);
    
    HIEFFPLA_INST_0_56592 : MX2
      port map(A => HIEFFPLA_NET_0_75201, B => 
        HIEFFPLA_NET_0_75075, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75234);
    
    HIEFFPLA_INST_0_65099 : AOI1D
      port map(A => HIEFFPLA_NET_0_73454, B => 
        HIEFFPLA_NET_0_73453, C => 
        \Pressure_Signal_Debounce_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73472);
    
    HIEFFPLA_INST_0_57887 : AO1B
      port map(A => \Sensors_0_pressure_time[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, C
         => HIEFFPLA_NET_0_74914, Y => HIEFFPLA_NET_0_74915);
    
    \General_Controller_0/uc_tx_state[1]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73572, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[1]_net_1\);
    
    HIEFFPLA_INST_0_67160 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[3]_net_1\, 
        B => HIEFFPLA_NET_0_72955, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72949);
    
    HIEFFPLA_INST_0_57044 : AOI1D
      port map(A => HIEFFPLA_NET_0_74839, B => 
        HIEFFPLA_NET_0_74951, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75177);
    
    HIEFFPLA_INST_0_69799 : NOR2A
      port map(A => HIEFFPLA_NET_0_72236, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72300);
    
    HIEFFPLA_INST_0_61224 : OR3B
      port map(A => 
        \General_Controller_0/state_seconds[13]_net_1\, B => 
        \General_Controller_0/state_seconds[12]_net_1\, C => 
        HIEFFPLA_NET_0_74251, Y => HIEFFPLA_NET_0_74244);
    
    HIEFFPLA_INST_0_88364 : AO1
      port map(A => HIEFFPLA_NET_0_88386, B => 
        HIEFFPLA_NET_0_75341, C => HIEFFPLA_NET_0_88387, Y => 
        HIEFFPLA_NET_0_89701);
    
    HIEFFPLA_INST_0_70405 : XOR2
      port map(A => HIEFFPLA_NET_0_72161, B => 
        \Timekeeper_0_microseconds[15]\, Y => 
        HIEFFPLA_NET_0_72145);
    
    HIEFFPLA_INST_0_63956 : MX2
      port map(A => HIEFFPLA_NET_0_73656, B => 
        HIEFFPLA_NET_0_73648, S => HIEFFPLA_NET_0_73599, Y => 
        HIEFFPLA_NET_0_73685);
    
    HIEFFPLA_INST_0_65314 : AOI1B
      port map(A => HIEFFPLA_NET_0_73417, B => 
        HIEFFPLA_NET_0_73412, C => HIEFFPLA_NET_0_73277, Y => 
        HIEFFPLA_NET_0_73414);
    
    HIEFFPLA_INST_0_62717 : NAND3C
      port map(A => HIEFFPLA_NET_0_73884, B => 
        HIEFFPLA_NET_0_73889, C => HIEFFPLA_NET_0_73776, Y => 
        HIEFFPLA_NET_0_73922);
    
    HIEFFPLA_INST_0_66949 : NAND3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        B => HIEFFPLA_NET_0_72745, C => HIEFFPLA_NET_0_72998, Y
         => HIEFFPLA_NET_0_72999);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1E1C0_data_out[6]\\\\/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75281, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \FMC_DA_c[6]\);
    
    HIEFFPLA_INST_0_66869 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_we\, 
        C => HIEFFPLA_NET_0_73012, Y => HIEFFPLA_NET_0_73016);
    
    HIEFFPLA_INST_0_62794 : AO1
      port map(A => HIEFFPLA_NET_0_73800, B => 
        \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        HIEFFPLA_NET_0_73964, Y => HIEFFPLA_NET_0_73902);
    
    HIEFFPLA_INST_0_60899 : AND2B
      port map(A => 
        \General_Controller_0/constant_bias_probe_id[0]_net_1\, B
         => \General_Controller_0/un10_uc_tx_rdy_i[1]\, Y => 
        HIEFFPLA_NET_0_74325);
    
    HIEFFPLA_INST_0_55957 : NAND2B
      port map(A => HIEFFPLA_NET_0_75382, B => 
        HIEFFPLA_NET_0_75396, Y => HIEFFPLA_NET_0_75384);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[2]\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_73128, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73041, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[2]_net_1\);
    
    HIEFFPLA_INST_0_57700 : AOI1
      port map(A => \Sensors_0_mag_y[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_74965, Y => HIEFFPLA_NET_0_74966);
    
    HIEFFPLA_INST_0_59698 : MX2
      port map(A => HIEFFPLA_NET_0_74539, B => 
        HIEFFPLA_NET_0_74518, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74520);
    
    \GS_Readout_0/subState[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74352, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/subState[3]_net_1\);
    
    HIEFFPLA_INST_0_68914 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, B
         => \Sensors_0/Gyro_0/I2C_Master_0_s_ack_error\, C => 
        \Sensors_0/Gyro_0/state[8]\, Y => HIEFFPLA_NET_0_72523);
    
    \EMU_RX_pad/U0/U0\ : IOPAD_IN
      port map(PAD => EMU_RX, Y => \EMU_RX_pad/U0/NET1\);
    
    HIEFFPLA_INST_0_68283 : NAND3C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[2]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[1]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_72690);
    
    \Science_0/ADC_READ_0/chan3_data[9]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[9]\);
    
    HIEFFPLA_INST_0_57303 : AND2
      port map(A => \Sensors_0_gyro_time[21]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75082);
    
    HIEFFPLA_INST_0_69190 : AO1A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        B => HIEFFPLA_NET_0_72437, C => HIEFFPLA_NET_0_72450, Y
         => HIEFFPLA_NET_0_72451);
    
    HIEFFPLA_INST_0_57897 : AO1B
      port map(A => \Sensors_0_mag_time[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74911, Y => HIEFFPLA_NET_0_74912);
    
    HIEFFPLA_INST_0_64541 : AO1A
      port map(A => HIEFFPLA_NET_0_73562, B => 
        HIEFFPLA_NET_0_73611, C => HIEFFPLA_NET_0_73617, Y => 
        HIEFFPLA_NET_0_73604);
    
    \Science_0/ADC_READ_0/exp_packet_1[8]\ : DFN1E0
      port map(D => \AFLSDF_INV_22\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[8]\);
    
    \Science_0/ADC_RESET_0/state[1]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73232, CLK => \s_time[5]\, E
         => CLKINT_1_Y, Q => 
        \Science_0/ADC_RESET_0/state[1]_net_1\);
    
    AFLSDF_INV_28 : INV
      port map(A => Sensors_0_mag_new_data, Y => \AFLSDF_INV_28\);
    
    HIEFFPLA_INST_0_56778 : AOI1C
      port map(A => HIEFFPLA_NET_0_75174, B => 
        HIEFFPLA_NET_0_75175, C => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75211);
    
    HIEFFPLA_INST_0_62755 : AO1A
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => HIEFFPLA_NET_0_73950, C => HIEFFPLA_NET_0_73939, Y
         => HIEFFPLA_NET_0_73913);
    
    HIEFFPLA_INST_0_58137 : AO1
      port map(A => \Sensors_0_mag_time[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75149, Y => HIEFFPLA_NET_0_74842);
    
    HIEFFPLA_INST_0_55044 : AND3
      port map(A => HIEFFPLA_NET_0_75593, B => 
        HIEFFPLA_NET_0_75591, C => HIEFFPLA_NET_0_75564, Y => 
        HIEFFPLA_NET_0_75605);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[5]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[5]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[5]\);
    
    HIEFFPLA_INST_0_66976 : OA1C
      port map(A => HIEFFPLA_NET_0_72981, B => 
        HIEFFPLA_NET_0_72913, C => HIEFFPLA_NET_0_72992, Y => 
        HIEFFPLA_NET_0_72993);
    
    HIEFFPLA_INST_0_56672 : MX2
      port map(A => HIEFFPLA_NET_0_75193, B => 
        HIEFFPLA_NET_0_75056, S => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75226);
    
    HIEFFPLA_INST_0_56083 : NOR2A
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, B
         => HIEFFPLA_NET_0_75350, Y => HIEFFPLA_NET_0_75351);
    
    HIEFFPLA_INST_0_68400 : AO1
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, C => 
        \Sensors_0/Gyro_0/state[8]\, Y => HIEFFPLA_NET_0_72658);
    
    HIEFFPLA_INST_0_57288 : AND2
      port map(A => \Sensors_0_gyro_time[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75092);
    
    \General_Controller_0/st_waddr[4]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[4]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_waddr[4]\);
    
    \Timing_0/s_time[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72040, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_time[2]_net_1\);
    
    HIEFFPLA_INST_0_56406 : MX2
      port map(A => \FMC_DA_c[0]\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[0]\\\\\, S => 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\, Y => 
        HIEFFPLA_NET_0_75287);
    
    HIEFFPLA_INST_0_64688 : NOR3A
      port map(A => HIEFFPLA_NET_0_73611, B => 
        HIEFFPLA_NET_0_73562, C => HIEFFPLA_NET_0_73978, Y => 
        HIEFFPLA_NET_0_73564);
    
    HIEFFPLA_INST_0_63255 : AO1
      port map(A => HIEFFPLA_NET_0_73888, B => 
        HIEFFPLA_NET_0_73811, C => HIEFFPLA_NET_0_73787, Y => 
        HIEFFPLA_NET_0_73798);
    
    HIEFFPLA_INST_0_69205 : NOR3B
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, 
        B => HIEFFPLA_NET_0_72540, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        Y => HIEFFPLA_NET_0_72447);
    
    HIEFFPLA_INST_0_63105 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state_0[1]_net_1\, 
        B => HIEFFPLA_NET_0_73827, C => HIEFFPLA_NET_0_73809, Y
         => HIEFFPLA_NET_0_73828);
    
    HIEFFPLA_INST_0_66756 : NAND3C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_73044);
    
    HIEFFPLA_INST_0_57778 : AOI1
      port map(A => \Science_0_exp_packet_0[51]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74783, Y => HIEFFPLA_NET_0_74945);
    
    HIEFFPLA_INST_0_61573 : AND3C
      port map(A => HIEFFPLA_NET_0_74180, B => 
        \General_Controller_0/sweep_table_probe_id[6]_net_1\, C
         => \General_Controller_0/sweep_table_probe_id[7]_net_1\, 
        Y => HIEFFPLA_NET_0_74181);
    
    \Science_0/ADC_READ_0/data_b[10]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[10]_net_1\);
    
    HIEFFPLA_INST_0_68178 : NOR3A
      port map(A => HIEFFPLA_NET_0_72772, B => 
        HIEFFPLA_NET_0_72902, C => HIEFFPLA_NET_0_72764, Y => 
        HIEFFPLA_NET_0_72714);
    
    \Eject_Signal_Debounce_0/ffu_ejected_out\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74751, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72220, Q => 
        Eject_Signal_Debounce_0_ffu_ejected_out);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[12]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72283, Q => 
        \Sensors_0_pressure_temp_raw[12]\);
    
    HIEFFPLA_INST_0_70502 : AX1C
      port map(A => \Timekeeper_0_milliseconds[17]\, B => 
        HIEFFPLA_NET_0_72121, C => 
        \Timekeeper_0_milliseconds[18]\, Y => 
        HIEFFPLA_NET_0_72107);
    
    HIEFFPLA_INST_0_60056 : AND2B
      port map(A => HIEFFPLA_NET_0_74371, B => 
        HIEFFPLA_NET_0_74552, Y => HIEFFPLA_NET_0_74468);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72465, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]_net_1\);
    
    HIEFFPLA_INST_0_69933 : AO1
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[3]_net_1\, 
        B => HIEFFPLA_NET_0_72238, C => HIEFFPLA_NET_0_72258, Y
         => HIEFFPLA_NET_0_72264);
    
    HIEFFPLA_INST_0_57762 : AOI1
      port map(A => \Science_0_exp_packet_0[62]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74814, Y => HIEFFPLA_NET_0_74950);
    
    HIEFFPLA_INST_0_69290 : NOR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72428);
    
    HIEFFPLA_INST_0_67450 : OR2A
      port map(A => HIEFFPLA_NET_0_72875, B => 
        HIEFFPLA_NET_0_72764, Y => HIEFFPLA_NET_0_72876);
    
    \Science_0/ADC_READ_0/exp_packet_1[46]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[12]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[46]\);
    
    HIEFFPLA_INST_0_70487 : XOR2
      port map(A => HIEFFPLA_NET_0_72119, B => 
        \Timekeeper_0_milliseconds[11]\, Y => 
        HIEFFPLA_NET_0_72114);
    
    HIEFFPLA_INST_0_64612 : AND2B
      port map(A => \General_Controller_0/uc_tx_state[5]_net_1\, 
        B => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73587);
    
    HIEFFPLA_INST_0_61769 : XOR2
      port map(A => HIEFFPLA_NET_0_74147, B => 
        \General_Controller_0/sweep_table_sweep_cnt[13]_net_1\, Y
         => HIEFFPLA_NET_0_74140);
    
    HIEFFPLA_INST_0_55167 : NOR3A
      port map(A => HIEFFPLA_NET_0_75579, B => 
        HIEFFPLA_NET_0_75567, C => HIEFFPLA_NET_0_75578, Y => 
        HIEFFPLA_NET_0_75570);
    
    HIEFFPLA_INST_0_69450 : AO1
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        B => PRESSURE_SCL_c, C => HIEFFPLA_NET_0_72347, Y => 
        HIEFFPLA_NET_0_72385);
    
    \General_Controller_0/state_seconds[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74226, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[2]_net_1\);
    
    HIEFFPLA_INST_0_68527 : AO1A
      port map(A => GYRO_SCL_c, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, C => 
        CLKINT_1_Y, Y => HIEFFPLA_NET_0_72627);
    
    HIEFFPLA_INST_0_61404 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[43]\, B => 
        \Timekeeper_0_milliseconds[3]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74203);
    
    \General_Controller_0/status_bits_1[59]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74187, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[59]\);
    
    HIEFFPLA_INST_0_60367 : AND2B
      port map(A => HIEFFPLA_NET_0_74556, B => 
        HIEFFPLA_NET_0_74459, Y => HIEFFPLA_NET_0_74426);
    
    HIEFFPLA_INST_0_61639 : MX2
      port map(A => \SweepTable_0_RD[11]\, B => 
        \SweepTable_1_RD[11]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74168);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[3]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72503, Q => 
        \Sensors_0_gyro_x[3]\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/data_out[3]\ : DFN0E1C1
      port map(D => GYRO_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72680, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[5]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72783, Q => 
        \Sensors_0_mag_y[5]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[4]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72215, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[4]_net_1\);
    
    HIEFFPLA_INST_0_66221 : XOR2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G2[1]_net_1\, B
         => \Science_0/ADC_READ_0_G2[1]\, Y => 
        HIEFFPLA_NET_0_73174);
    
    \PRESSURE_SCL_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => PRESSURE_SCL_c, E => \VCC\, DOUT => 
        \PRESSURE_SCL_pad/U0/NET1\, EOUT => 
        \PRESSURE_SCL_pad/U0/NET2\);
    
    \Timing_0/f_time[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72087, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/f_time[3]_net_1\);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[5]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_75248, CLK => CLKINT_0_Y_0, E
         => CLKINT_1_Y, Q => 
        \Data_Saving_0/Interrupt_Generator_0/counter[5]_net_1\);
    
    HIEFFPLA_INST_0_70769 : AO1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_s_ack_error\, B
         => HIEFFPLA_NET_0_72015, C => HIEFFPLA_NET_0_72259, Y
         => HIEFFPLA_NET_0_72265);
    
    HIEFFPLA_INST_0_61160 : AOI1C
      port map(A => HIEFFPLA_NET_0_74245, B => 
        HIEFFPLA_NET_0_74247, C => 
        \General_Controller_0/state_seconds[7]_net_1\, Y => 
        HIEFFPLA_NET_0_74260);
    
    HIEFFPLA_INST_0_58381 : AND2
      port map(A => \Sensors_0_mag_z[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        Y => HIEFFPLA_NET_0_74785);
    
    \GS_Readout_0/state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74614, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/state[0]_net_1\);
    
    HIEFFPLA_INST_0_67387 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, C
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72895);
    
    HIEFFPLA_INST_0_64968 : OR3A
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[7]_net_1\, 
        B => \Pressure_Signal_Debounce_0/ms_cnt[4]_net_1\, C => 
        \Pressure_Signal_Debounce_0/ms_cnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73500);
    
    \Communications_0/UART_1/tx_clk_count[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75411, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_clk_count[0]_net_1\);
    
    HIEFFPLA_INST_0_60843 : AND2
      port map(A => HIEFFPLA_NET_0_74345, B => 
        \GS_Readout_0/subState[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74346);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRYSYNC[2]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_5_Q\, CLK
         => CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[2]\\\\\);
    
    HIEFFPLA_INST_0_58382 : AND2
      port map(A => \Sensors_0_mag_z[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        Y => HIEFFPLA_NET_0_74784);
    
    HIEFFPLA_INST_0_58087 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[13]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75154, Y => HIEFFPLA_NET_0_74858);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[9]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72782, Q => 
        \Sensors_0_mag_y[9]\);
    
    HIEFFPLA_INST_0_55130 : NOR3B
      port map(A => HIEFFPLA_NET_0_75596, B => 
        \Communications_0/UART_0/rx_clk_count[24]_net_1\, C => 
        \Communications_0/UART_0/rx_clk_count[23]_net_1\, Y => 
        HIEFFPLA_NET_0_75581);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73037, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\);
    
    HIEFFPLA_INST_0_56889 : MX2
      port map(A => HIEFFPLA_NET_0_74996, B => 
        HIEFFPLA_NET_0_74924, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75199);
    
    HIEFFPLA_INST_0_56464 : XNOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[4]\\\\\, B => 
        HIEFFPLA_NET_0_75273, Y => HIEFFPLA_NET_0_75274);
    
    \FMC_DA_pad[6]/U0/U1\ : IOTRI_OB_EB
      port map(D => \FMC_DA_c[6]\, E => \VCC\, DOUT => 
        \FMC_DA_pad[6]/U0/NET1\, EOUT => \FMC_DA_pad[6]/U0/NET2\);
    
    \Science_0/ADC_READ_0/chan2_data[7]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[7]\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRY[5]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75309, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[5]\\\\\);
    
    HIEFFPLA_INST_0_61288 : XA1B
      port map(A => \General_Controller_0/state_seconds[0]_net_1\, 
        B => \General_Controller_0/state_seconds[1]_net_1\, C => 
        HIEFFPLA_NET_0_74217, Y => HIEFFPLA_NET_0_74227);
    
    HIEFFPLA_INST_0_55437 : NOR3A
      port map(A => 
        \Communications_0/UART_0/tx_clk_count[1]_net_1\, B => 
        \Communications_0/UART_0/tx_state[0]_net_1\, C => 
        \Communications_0/UART_0/tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75513);
    
    HIEFFPLA_INST_0_62907 : AO1
      port map(A => HIEFFPLA_NET_0_73861, B => 
        HIEFFPLA_NET_0_73775, C => HIEFFPLA_NET_0_74075, Y => 
        HIEFFPLA_NET_0_73868);
    
    \Timekeeper_0/milliseconds[20]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72104, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[20]\);
    
    HIEFFPLA_INST_0_67397 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        C => HIEFFPLA_NET_0_72761, Y => HIEFFPLA_NET_0_72892);
    
    HIEFFPLA_INST_0_67087 : NOR2A
      port map(A => HIEFFPLA_NET_0_72963, B => 
        HIEFFPLA_NET_0_72964, Y => HIEFFPLA_NET_0_72967);
    
    HIEFFPLA_INST_0_68524 : AO1A
      port map(A => GYRO_SDA_in, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, C => 
        HIEFFPLA_NET_0_72627, Y => HIEFFPLA_NET_0_72628);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[13]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[13]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[13]\);
    
    HIEFFPLA_INST_0_60033 : MX2
      port map(A => \Sensors_0_pressure_raw[17]\, B => 
        \Sensors_0_pressure_raw[21]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74471);
    
    HIEFFPLA_INST_0_56442 : MX2
      port map(A => \FMC_DA_c[6]\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[6]\\\\\, S => 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\, Y => 
        HIEFFPLA_NET_0_75281);
    
    HIEFFPLA_INST_0_62801 : OA1A
      port map(A => HIEFFPLA_NET_0_73897, B => 
        HIEFFPLA_NET_0_73988, C => HIEFFPLA_NET_0_73937, Y => 
        HIEFFPLA_NET_0_73899);
    
    HIEFFPLA_INST_0_55133 : NAND3
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[29]_net_1\, B => 
        \Communications_0/UART_0/rx_clk_count_c0\, C => 
        \Communications_0/UART_0/rx_clk_count[30]_net_1\, Y => 
        HIEFFPLA_NET_0_75579);
    
    HIEFFPLA_INST_0_57420 : AO1
      port map(A => \Science_0_exp_packet_0[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74849, Y => HIEFFPLA_NET_0_75051);
    
    HIEFFPLA_INST_0_67794 : AND3C
      port map(A => HIEFFPLA_NET_0_72765, B => 
        HIEFFPLA_NET_0_72900, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72800);
    
    HIEFFPLA_INST_0_64786 : AO1
      port map(A => Communications_0_uc_tx_rdy, B => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, C => 
        \General_Controller_0/uc_tx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73541);
    
    HIEFFPLA_INST_0_60308 : MX2
      port map(A => HIEFFPLA_NET_0_74385, B => 
        HIEFFPLA_NET_0_74358, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74433);
    
    HIEFFPLA_INST_0_68796 : AND2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, B
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        Y => HIEFFPLA_NET_0_72558);
    
    \General_Controller_0/constant_bias_probe_id[3]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73923, Q => 
        \General_Controller_0/un10_uc_tx_rdy_i[3]\);
    
    HIEFFPLA_INST_0_57927 : AO1B
      port map(A => \Sensors_0_mag_time[12]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74902, Y => HIEFFPLA_NET_0_74903);
    
    HIEFFPLA_INST_0_58567 : NOR3B
      port map(A => \Eject_Signal_Debounce_0/ms_cnt[0]_net_1\, B
         => HIEFFPLA_NET_0_74737, C => HIEFFPLA_NET_0_74739, Y
         => HIEFFPLA_NET_0_74733);
    
    HIEFFPLA_INST_0_65155 : AOI1C
      port map(A => HIEFFPLA_NET_0_73459, B => 
        HIEFFPLA_NET_0_73462, C => \Sensors_0_pressure_raw[19]\, 
        Y => HIEFFPLA_NET_0_73456);
    
    HIEFFPLA_INST_0_64611 : AND2B
      port map(A => \General_Controller_0/uc_tx_state[3]_net_1\, 
        B => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73588);
    
    HIEFFPLA_INST_0_65279 : NAND2B
      port map(A => \Science_0/ADC_READ_0/state[2]_net_1\, B => 
        \Science_0/ADC_READ_0/countere\, Y => 
        HIEFFPLA_NET_0_73425);
    
    HIEFFPLA_INST_0_59073 : NAND2B
      port map(A => HIEFFPLA_NET_0_74633, B => 
        HIEFFPLA_NET_0_74620, Y => HIEFFPLA_NET_0_74621);
    
    HIEFFPLA_INST_0_65108 : AND3B
      port map(A => HIEFFPLA_NET_0_73467, B => 
        HIEFFPLA_NET_0_73459, C => 
        \Pressure_Signal_Debounce_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73470);
    
    HIEFFPLA_INST_0_62274 : OA1A
      port map(A => HIEFFPLA_NET_0_73948, B => 
        HIEFFPLA_NET_0_74072, C => HIEFFPLA_NET_0_74034, Y => 
        HIEFFPLA_NET_0_74016);
    
    \General_Controller_0/temp_first_byte[1]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73872, Q => 
        \General_Controller_0/temp_first_byte[1]_net_1\);
    
    \General_Controller_0/st_raddr[1]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[1]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73979, Q => 
        \General_Controller_0_st_raddr_1[1]\);
    
    HIEFFPLA_INST_0_62307 : AO1A
      port map(A => HIEFFPLA_NET_0_73914, B => 
        \General_Controller_0/uc_rx_state[0]_net_1\, C => 
        HIEFFPLA_NET_0_73874, Y => HIEFFPLA_NET_0_74009);
    
    HIEFFPLA_INST_0_60699 : MX2
      port map(A => \Science_0_chan2_data[6]\, B => 
        \Science_0_chan2_data[10]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74375);
    
    HIEFFPLA_INST_0_67585 : NOR3A
      port map(A => HIEFFPLA_NET_0_72839, B => 
        HIEFFPLA_NET_0_72929, C => HIEFFPLA_NET_0_72935, Y => 
        HIEFFPLA_NET_0_72847);
    
    HIEFFPLA_INST_0_55186 : AX1A
      port map(A => HIEFFPLA_NET_0_75579, B => 
        \Communications_0/UART_0/rx_clk_count[28]_net_1\, C => 
        \Communications_0/UART_0/rx_clk_count[27]_net_1\, Y => 
        HIEFFPLA_NET_0_75565);
    
    HIEFFPLA_INST_0_61754 : AND3
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[7]_net_1\, B
         => HIEFFPLA_NET_0_74145, C => 
        \General_Controller_0/sweep_table_sweep_cnt[8]_net_1\, Y
         => HIEFFPLA_NET_0_74146);
    
    HIEFFPLA_INST_0_57707 : AO1B
      port map(A => \Sensors_0_pressure_raw[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74963, Y => HIEFFPLA_NET_0_74964);
    
    HIEFFPLA_INST_0_67090 : NAND2B
      port map(A => HIEFFPLA_NET_0_72964, B => 
        HIEFFPLA_NET_0_72962, Y => HIEFFPLA_NET_0_72966);
    
    \Data_Saving_0/Packet_Saver_0/old_ch_0_new_data\ : DFN0P1
      port map(D => \AFLSDF_INV_23\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => 
        \Data_Saving_0/Packet_Saver_0/old_ch_0_new_data_i_0\);
    
    HIEFFPLA_INST_0_71005 : OR3B
      port map(A => \Pressure_Signal_Debounce_0/state[1]_net_1\, 
        B => \Sensors_0_pressure_raw[22]\, C => 
        HIEFFPLA_NET_0_73471, Y => HIEFFPLA_NET_0_71993);
    
    \General_Controller_0/st_raddr[3]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[3]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73979, Q => 
        \General_Controller_0_st_raddr_1[3]\);
    
    \LDCLK_pad/U0/U0\ : IOPAD_TRI
      port map(D => \LDCLK_pad/U0/NET1\, E => \LDCLK_pad/U0/NET2\, 
        PAD => LDCLK);
    
    HIEFFPLA_INST_0_57690 : AOI1
      port map(A => \Sensors_0_acc_y[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74968, Y => HIEFFPLA_NET_0_74969);
    
    HIEFFPLA_INST_0_55256 : NOR3B
      port map(A => HIEFFPLA_NET_0_75550, B => 
        \Communications_0/UART_0/rx_state[0]_net_1\, C => 
        HIEFFPLA_NET_0_75582, Y => HIEFFPLA_NET_0_75551);
    
    HIEFFPLA_INST_0_55433 : AX1B
      port map(A => HIEFFPLA_NET_0_75536, B => 
        \Communications_0/UART_0/tx_clk_count_i_0[3]\, C => 
        \Communications_0/UART_0/tx_clk_count_i_0[4]\, Y => 
        HIEFFPLA_NET_0_75514);
    
    \Timing_0/m_time[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72065, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \s_clks_net_0[9]\);
    
    HIEFFPLA_INST_0_61786 : XOR2
      port map(A => HIEFFPLA_NET_0_74150, B => 
        \General_Controller_0/sweep_table_sweep_cnt[5]_net_1\, Y
         => HIEFFPLA_NET_0_74133);
    
    \General_Controller_0/sweep_table_sweep_cnt[8]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74130, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[8]_net_1\);
    
    HIEFFPLA_INST_0_66114 : AOI1A
      port map(A => \Science_0/DAC_SET_0/old_set_net_1\, B => 
        \Science_0/SWEEP_SPIDER2_0_SET\, C => LDCLK_c, Y => 
        HIEFFPLA_NET_0_73206);
    
    HIEFFPLA_INST_0_61233 : OR3B
      port map(A => \General_Controller_0/state_seconds[8]_net_1\, 
        B => \General_Controller_0/state_seconds[9]_net_1\, C => 
        HIEFFPLA_NET_0_74261, Y => HIEFFPLA_NET_0_74241);
    
    HIEFFPLA_INST_0_57141 : AND2
      port map(A => \Sensors_0_pressure_temp_raw[21]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75156);
    
    HIEFFPLA_INST_0_55050 : AND3C
      port map(A => \Communications_0/UART_0/rx_count[2]_net_1\, 
        B => \Communications_0/UART_0/rx_count[1]_net_1\, C => 
        \Communications_0/UART_0/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75603);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[1]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72767, Q => 
        \Sensors_0_acc_y[1]\);
    
    HIEFFPLA_INST_0_66771 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        B => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73038);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[20]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72280, Q => \Sensors_0_pressure_raw[20]\);
    
    HIEFFPLA_INST_0_59991 : MX2
      port map(A => \Science_0_chan3_data[1]\, B => 
        \Science_0_chan3_data[5]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74477);
    
    HIEFFPLA_INST_0_65257 : NOR3A
      port map(A => HIEFFPLA_NET_0_73432, B => 
        \Sensors_0_pressure_raw[15]\, C => 
        \Sensors_0_pressure_raw[17]\, Y => HIEFFPLA_NET_0_73433);
    
    \General_Controller_0/state_seconds[10]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74239, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[10]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[14]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72553, Q => 
        \Sensors_0_gyro_x[14]\);
    
    HIEFFPLA_INST_0_56510 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, B
         => HIEFFPLA_NET_0_75349, Y => HIEFFPLA_NET_0_75259);
    
    HIEFFPLA_INST_0_68906 : NOR3B
      port map(A => HIEFFPLA_NET_0_72508, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72525);
    
    HIEFFPLA_INST_0_71117 : AOI1D
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => \Sensors_0_acc_temp[1]\, Y => HIEFFPLA_NET_0_71980);
    
    HIEFFPLA_INST_0_62007 : AND3
      port map(A => HIEFFPLA_NET_0_74113, B => 
        HIEFFPLA_NET_0_74111, C => HIEFFPLA_NET_0_74092, Y => 
        HIEFFPLA_NET_0_74075);
    
    HIEFFPLA_INST_0_58125 : AO1
      port map(A => \Sensors_0_mag_time[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75152, Y => HIEFFPLA_NET_0_74845);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[15]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72281, Q => \Sensors_0_pressure_raw[15]\);
    
    HIEFFPLA_INST_0_65520 : AND2
      port map(A => \Science_0/ADC_READ_0/cnt3dn[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt3dn[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73354);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[7]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75260, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[7]\\\\\);
    
    HIEFFPLA_INST_0_62000 : AND2B
      port map(A => \General_Controller_0/uc_rx_byte[7]_net_1\, B
         => \General_Controller_0/uc_rx_byte[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74077);
    
    HIEFFPLA_INST_0_68528 : NOR2A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, B => 
        GYRO_SCL_c, Y => HIEFFPLA_NET_0_72626);
    
    HIEFFPLA_INST_0_61699 : MX2
      port map(A => \SweepTable_0_RD[6]\, B => 
        \SweepTable_1_RD[6]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74158);
    
    HIEFFPLA_INST_0_65428 : OR2A
      port map(A => \Science_0/ADC_READ_0/cnt2dn[4]_net_1\, B => 
        HIEFFPLA_NET_0_73387, Y => HIEFFPLA_NET_0_73379);
    
    HIEFFPLA_INST_0_71128 : AO1
      port map(A => \Science_0_exp_packet_0[36]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74835, Y => HIEFFPLA_NET_0_71978);
    
    HIEFFPLA_INST_0_68644 : AO1A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_we\, C => 
        HIEFFPLA_NET_0_72588, Y => HIEFFPLA_NET_0_72598);
    
    HIEFFPLA_INST_0_57515 : AO1
      port map(A => \Sensors_0_acc_z[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74858, Y => HIEFFPLA_NET_0_75023);
    
    HIEFFPLA_INST_0_65809 : NOR3A
      port map(A => HIEFFPLA_NET_0_73275, B => 
        \Science_0/ADC_READ_0/data_b[17]_net_1\, C => 
        \Science_0/ADC_READ_0/data_b[16]_net_1\, Y => 
        HIEFFPLA_NET_0_73276);
    
    HIEFFPLA_INST_0_65637 : NOR3A
      port map(A => \Science_0/ADC_READ_0/cnt4dn[3]_net_1\, B => 
        HIEFFPLA_NET_0_73320, C => 
        \Science_0/ADC_READ_0/cnt4dn[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73321);
    
    HIEFFPLA_INST_0_56905 : MX2
      port map(A => HIEFFPLA_NET_0_74990, B => 
        HIEFFPLA_NET_0_74918, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75197);
    
    HIEFFPLA_INST_0_69240 : AO1A
      port map(A => HIEFFPLA_NET_0_72479, B => 
        HIEFFPLA_NET_0_72551, C => HIEFFPLA_NET_0_72440, Y => 
        HIEFFPLA_NET_0_72441);
    
    HIEFFPLA_INST_0_63089 : NOR3B
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, C => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73832);
    
    HIEFFPLA_INST_0_60720 : MX2
      port map(A => HIEFFPLA_NET_0_74480, B => 
        HIEFFPLA_NET_0_74417, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74370);
    
    \Timing_0/m_count[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72027, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_count[1]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[6]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72489, Q => 
        \ch3_data_net_0[2]\);
    
    HIEFFPLA_INST_0_63590 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[9]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_sample_skip[9]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73744);
    
    HIEFFPLA_INST_0_62881 : AO1
      port map(A => HIEFFPLA_NET_0_73800, B => 
        \General_Controller_0/uc_rx_state[3]_net_1\, C => 
        HIEFFPLA_NET_0_73962, Y => HIEFFPLA_NET_0_73876);
    
    HIEFFPLA_INST_0_68756 : AOI1
      port map(A => HIEFFPLA_NET_0_72506, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, C
         => HIEFFPLA_NET_0_72566, Y => HIEFFPLA_NET_0_72569);
    
    HIEFFPLA_INST_0_67134 : NOR3A
      port map(A => HIEFFPLA_NET_0_72879, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[8]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72957);
    
    HIEFFPLA_INST_0_61948 : NOR3B
      port map(A => HIEFFPLA_NET_0_73907, B => 
        HIEFFPLA_NET_0_74074, C => HIEFFPLA_NET_0_73810, Y => 
        HIEFFPLA_NET_0_74091);
    
    HIEFFPLA_INST_0_59025 : OA1A
      port map(A => HIEFFPLA_NET_0_74405, B => 
        HIEFFPLA_NET_0_74500, C => \GS_Readout_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_74633);
    
    HIEFFPLA_INST_0_56507 : AX1C
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, B
         => HIEFFPLA_NET_0_75352, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[7]\\\\\, Y
         => HIEFFPLA_NET_0_75260);
    
    HIEFFPLA_INST_0_62597 : AND3B
      port map(A => 
        \General_Controller_0/uc_rx_substate[4]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[3]_net_1\, C => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73949);
    
    \Science_0/ADC_READ_0/data_b[9]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[9]_net_1\);
    
    HIEFFPLA_INST_0_55141 : XA1B
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[23]_net_1\, B => 
        HIEFFPLA_NET_0_75566, C => HIEFFPLA_NET_0_75567, Y => 
        HIEFFPLA_NET_0_75576);
    
    \General_Controller_0/sweep_table_sample_skip[13]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[13]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[14]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[14]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[14]\);
    
    HIEFFPLA_INST_0_62552 : OR3A
      port map(A => HIEFFPLA_NET_0_73897, B => 
        HIEFFPLA_NET_0_73882, C => HIEFFPLA_NET_0_73988, Y => 
        HIEFFPLA_NET_0_73958);
    
    HIEFFPLA_INST_0_69812 : XA1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[3]_net_1\, 
        B => HIEFFPLA_NET_0_72307, C => HIEFFPLA_NET_0_72236, Y
         => HIEFFPLA_NET_0_72297);
    
    HIEFFPLA_INST_0_58504 : OA1C
      port map(A => HIEFFPLA_NET_0_74738, B => 
        HIEFFPLA_NET_0_74732, C => HIEFFPLA_NET_0_74740, Y => 
        HIEFFPLA_NET_0_74747);
    
    HIEFFPLA_INST_0_69956 : AOI1D
      port map(A => HIEFFPLA_NET_0_72228, B => 
        HIEFFPLA_NET_0_72243, C => HIEFFPLA_NET_0_72254, Y => 
        HIEFFPLA_NET_0_72260);
    
    HIEFFPLA_INST_0_65755 : XA1B
      port map(A => HIEFFPLA_NET_0_73297, B => 
        \Science_0/ADC_READ_0/cnt[3]_net_1\, C => 
        HIEFFPLA_NET_0_73241, Y => HIEFFPLA_NET_0_73288);
    
    \Science_0/ADC_READ_0/exp_packet_1[44]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[10]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[44]\);
    
    HIEFFPLA_INST_0_56012 : AND3A
      port map(A => \Data_Saving_0/FPGA_Buffer_0/empty\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[0]\\\\\, C
         => FMC_NOE_c, Y => HIEFFPLA_NET_0_75369);
    
    \General_Controller_0/st_raddr[0]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[0]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73979, Q => 
        \General_Controller_0_st_raddr_1[0]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[38]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[4]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[38]\);
    
    HIEFFPLA_INST_0_67466 : AND3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        C => HIEFFPLA_NET_0_72871, Y => HIEFFPLA_NET_0_72872);
    
    \ARST_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => ARST_c, E => \VCC\, DOUT => 
        \ARST_pad/U0/NET1\, EOUT => \ARST_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_67346 : AND3A
      port map(A => \Sensors_0/Accelerometer_0/state[8]\, B => 
        HIEFFPLA_NET_0_72759, C => HIEFFPLA_NET_0_72929, Y => 
        HIEFFPLA_NET_0_72902);
    
    HIEFFPLA_INST_0_66666 : AND3C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        C => \Sensors_0/Accelerometer_0/state_0[8]\, Y => 
        HIEFFPLA_NET_0_73070);
    
    \General_Controller_0/sweep_table_samples_per_step[10]\ : 
        DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[2]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[10]_net_1\);
    
    HIEFFPLA_INST_0_67507 : NAND3C
      port map(A => HIEFFPLA_NET_0_72850, B => 
        HIEFFPLA_NET_0_72860, C => HIEFFPLA_NET_0_72861, Y => 
        HIEFFPLA_NET_0_72862);
    
    HIEFFPLA_INST_0_64417 : MX2
      port map(A => HIEFFPLA_NET_0_73708, B => 
        HIEFFPLA_NET_0_73700, S => HIEFFPLA_NET_0_73593, Y => 
        HIEFFPLA_NET_0_73628);
    
    HIEFFPLA_INST_0_57340 : AO1B
      port map(A => \Sensors_0_pressure_temp_raw[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_75071, Y => HIEFFPLA_NET_0_75072);
    
    HIEFFPLA_INST_0_70663 : XA1B
      port map(A => \Timing_0/s_count[6]_net_1\, B => 
        HIEFFPLA_NET_0_72019, C => HIEFFPLA_NET_0_72058, Y => 
        HIEFFPLA_NET_0_72051);
    
    HIEFFPLA_INST_0_69978 : NOR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_s_ack_error\, Y
         => HIEFFPLA_NET_0_72254);
    
    HIEFFPLA_INST_0_68943 : NAND3
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, C
         => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, Y => 
        HIEFFPLA_NET_0_72516);
    
    HIEFFPLA_INST_0_57468 : AOI1
      port map(A => \Science_0_exp_packet_0[29]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_75036, Y => HIEFFPLA_NET_0_75037);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_WADDR[0]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75331, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[0]\\\\\);
    
    HIEFFPLA_INST_0_70408 : AX1C
      port map(A => \Timekeeper_0_microseconds[15]\, B => 
        HIEFFPLA_NET_0_72161, C => 
        \Timekeeper_0_microseconds[16]\, Y => 
        HIEFFPLA_NET_0_72144);
    
    HIEFFPLA_INST_0_70397 : XOR2
      port map(A => HIEFFPLA_NET_0_72152, B => 
        \Timekeeper_0_microseconds[11]\, Y => 
        HIEFFPLA_NET_0_72149);
    
    HIEFFPLA_INST_0_69298 : NOR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\, 
        B => HIEFFPLA_NET_0_72345, C => HIEFFPLA_NET_0_72427, Y
         => HIEFFPLA_NET_0_72425);
    
    HIEFFPLA_INST_0_63536 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[8]_net_1\, B
         => \General_Controller_0/sweep_table_points[8]_net_1\, S
         => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73753);
    
    \General_Controller_0/sweep_table_read_value[4]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74160, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[4]_net_1\);
    
    HIEFFPLA_INST_0_70443 : AND3
      port map(A => \Timekeeper_0_milliseconds[11]\, B => 
        HIEFFPLA_NET_0_72119, C => 
        \Timekeeper_0_milliseconds[12]\, Y => 
        HIEFFPLA_NET_0_72127);
    
    HIEFFPLA_INST_0_55914 : AND2
      port map(A => HIEFFPLA_NET_0_75395, B => 
        \Communications_0/UART_1/tx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75396);
    
    HIEFFPLA_INST_0_62087 : AO1C
      port map(A => HIEFFPLA_NET_0_73875, B => 
        \General_Controller_0/uc_rx_prev_state[3]_net_1\, C => 
        HIEFFPLA_NET_0_73890, Y => HIEFFPLA_NET_0_74055);
    
    HIEFFPLA_INST_0_58378 : AND2
      port map(A => \Sensors_0_mag_z[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        Y => HIEFFPLA_NET_0_74786);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[7]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[7]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[7]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[3]\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72297, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72221, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[3]_net_1\);
    
    HIEFFPLA_INST_0_70537 : XOR2
      port map(A => \Timing_0/f_time[1]_net_1\, B => 
        \Timing_0/f_time[0]_net_1\, Y => HIEFFPLA_NET_0_72089);
    
    HIEFFPLA_INST_0_66993 : NAND3C
      port map(A => HIEFFPLA_NET_0_72987, B => 
        HIEFFPLA_NET_0_72983, C => HIEFFPLA_NET_0_72979, Y => 
        HIEFFPLA_NET_0_72988);
    
    HIEFFPLA_INST_0_60811 : AX1
      port map(A => Communications_0_ext_tx_rdy, B => 
        \GS_Readout_0/state[6]_net_1\, C => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74355);
    
    HIEFFPLA_INST_0_70973 : ZOR3I
      port map(A => \Science_0/ADC_READ_0/data_b[14]_net_1\, B
         => \Science_0/ADC_READ_0/data_b[13]_net_1\, C => 
        \Science_0/ADC_READ_0/data_b[12]_net_1\, Y => 
        HIEFFPLA_NET_0_71997);
    
    HIEFFPLA_INST_0_57880 : AOI1
      port map(A => \Sensors_0_acc_time[23]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74916, Y => HIEFFPLA_NET_0_74917);
    
    \General_Controller_0/uc_rx_prev_state[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74056, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_prev_state[2]_net_1\);
    
    \Science_0/ADC_READ_0/chan1_data[1]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[1]\);
    
    HIEFFPLA_INST_0_65510 : AX1C
      port map(A => \Science_0/ADC_READ_0/cnt2up[0]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2up[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt2up[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73359);
    
    \Science_0/ADC_READ_0/data_a[14]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[14]_net_1\);
    
    HIEFFPLA_INST_0_61012 : NOR2A
      port map(A => HIEFFPLA_NET_0_74294, B => 
        HIEFFPLA_NET_0_74259, Y => HIEFFPLA_NET_0_74295);
    
    \Science_0/ADC_READ_0/exp_packet_1[30]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[14]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[30]\);
    
    HIEFFPLA_INST_0_61335 : AX1C
      port map(A => \General_Controller_0/state_seconds[0]_net_1\, 
        B => \General_Controller_0/state_seconds[1]_net_1\, C => 
        \General_Controller_0/state_seconds[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74214);
    
    \FRAM_SCL_pad/U0/U0\ : IOPAD_TRI
      port map(D => \FRAM_SCL_pad/U0/NET1\, E => 
        \FRAM_SCL_pad/U0/NET2\, PAD => FRAM_SCL);
    
    HIEFFPLA_INST_0_55340 : MX2C
      port map(A => \Communications_0/UART_0/tx_byte[3]_net_1\, B
         => \Communications_0/UART_0/tx_byte[7]_net_1\, S => 
        \Communications_0/UART_0/tx_count[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75537);
    
    \Science_0/SET_LP_GAIN_0/old_G1[0]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73177, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/old_G1[0]_net_1\);
    
    HIEFFPLA_INST_0_65103 : OR3B
      port map(A => HIEFFPLA_NET_0_73470, B => 
        \Sensors_0_pressure_raw[20]\, C => HIEFFPLA_NET_0_73440, 
        Y => HIEFFPLA_NET_0_73471);
    
    \General_Controller_0/state_seconds[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74223, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[4]_net_1\);
    
    HIEFFPLA_INST_0_64950 : AND2B
      port map(A => \I2C_PassThrough_0.state[2]\, B => 
        \I2C_PassThrough_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73506);
    
    HIEFFPLA_INST_0_68614 : AOI1C
      port map(A => HIEFFPLA_NET_0_72599, B => 
        HIEFFPLA_NET_0_72585, C => HIEFFPLA_NET_0_72664, Y => 
        HIEFFPLA_NET_0_72605);
    
    HIEFFPLA_INST_0_67274 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72921);
    
    HIEFFPLA_INST_0_58490 : XNOR2
      port map(A => \Eject_Signal_Debounce_0/state[1]_net_1\, B
         => \Eject_Signal_Debounce_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74751);
    
    HIEFFPLA_INST_0_68361 : AO1A
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, C
         => HIEFFPLA_NET_0_72699, Y => HIEFFPLA_NET_0_72672);
    
    HIEFFPLA_INST_0_68041 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72747);
    
    \General_Controller_0/uc_rx_prev_state[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74054, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_prev_state[4]_net_1\);
    
    HIEFFPLA_INST_0_60434 : NOR2A
      port map(A => \Data_Hub_Packets_0_status_packet[3]\, B => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74415);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[4]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75263, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\);
    
    HIEFFPLA_INST_0_59020 : AND2B
      port map(A => \GS_Readout_0/state[3]_net_1\, B => 
        \GS_Readout_0/state[4]_net_1\, Y => HIEFFPLA_NET_0_74635);
    
    \Science_0/ADC_READ_0/chan5_data[0]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[0]\);
    
    HIEFFPLA_INST_0_64137 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_1[10]_net_1\, 
        B => 
        \General_Controller_0/constant_bias_voltage_1[2]_net_1\, 
        S => HIEFFPLA_NET_0_73558, Y => HIEFFPLA_NET_0_73663);
    
    HIEFFPLA_INST_0_57890 : AOI1
      port map(A => \Sensors_0_gyro_time[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74913, Y => HIEFFPLA_NET_0_74914);
    
    HIEFFPLA_INST_0_54987 : NAND3C
      port map(A => HIEFFPLA_NET_0_75618, B => 
        HIEFFPLA_NET_0_75617, C => HIEFFPLA_NET_0_75616, Y => 
        HIEFFPLA_NET_0_75619);
    
    \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_2\ : DFN0E0P1
      port map(D => HIEFFPLA_NET_0_72638, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72619, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_2_net_1\);
    
    \General_Controller_0/uc_tx_nextstate[1]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73625, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73857, Q => 
        \General_Controller_0/uc_tx_nextstate[1]_net_1\);
    
    \UC_I2C4_SDA_pad/U0/U1\ : IOBI_IB_OB_EB
      port map(D => \GND\, E => \I2C_PassThrough_0.state[2]\, YIN
         => \UC_I2C4_SDA_pad/U0/NET3\, DOUT => 
        \UC_I2C4_SDA_pad/U0/NET1\, EOUT => 
        \UC_I2C4_SDA_pad/U0/NET2\, Y => UC_I2C4_SDA_in);
    
    \Science_0/ADC_READ_0/cnt2up[2]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73362, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2up[2]_net_1\);
    
    HIEFFPLA_INST_0_69796 : AO1
      port map(A => HIEFFPLA_NET_0_72308, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[3]_net_1\, 
        C => HIEFFPLA_NET_0_72311, Y => HIEFFPLA_NET_0_72301);
    
    HIEFFPLA_INST_0_69780 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[2]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72308);
    
    HIEFFPLA_INST_0_55593 : AND2B
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[30]_net_1\, B => 
        \Communications_0/UART_1/rx_clk_count[29]_net_1\, Y => 
        HIEFFPLA_NET_0_75471);
    
    \General_Controller_0/unit_id[1]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73990, Q => 
        \General_Controller_0_unit_id[1]\);
    
    HIEFFPLA_INST_0_64691 : NAND3C
      port map(A => 
        \General_Controller_0/uc_tx_substate[0]_net_1\, B => 
        \General_Controller_0/uc_tx_substate[3]_net_1\, C => 
        \General_Controller_0/uc_tx_substate[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73563);
    
    \Science_0/ADC_READ_0/exp_packet_1[2]\ : DFN1E0
      port map(D => \AFLSDF_INV_24\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[2]\);
    
    HIEFFPLA_INST_0_60714 : NOR2A
      port map(A => HIEFFPLA_NET_0_74520, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74371);
    
    HIEFFPLA_INST_0_57226 : AO1
      port map(A => \Sensors_0_gyro_time[16]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75120, Y => HIEFFPLA_NET_0_75121);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[1]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72783, Q => 
        \Sensors_0_mag_y[1]\);
    
    HIEFFPLA_INST_0_55404 : XO1
      port map(A => HIEFFPLA_NET_0_75534, B => 
        \Communications_0/UART_0/tx_clk_count_i_0[6]\, C => 
        HIEFFPLA_NET_0_75527, Y => HIEFFPLA_NET_0_75520);
    
    HIEFFPLA_INST_0_57549 : AO1B
      port map(A => \Sensors_0_gyro_z[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75012, Y => HIEFFPLA_NET_0_75013);
    
    HIEFFPLA_INST_0_55138 : AND2
      port map(A => HIEFFPLA_NET_0_75586, B => 
        \Communications_0/UART_0/rx_clk_count[26]_net_1\, Y => 
        HIEFFPLA_NET_0_75577);
    
    \Science_0/ADC_READ_0/chan6_data[8]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[8]\);
    
    \Science_0/ADC_READ_0/chan0_data[8]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[8]\);
    
    HIEFFPLA_INST_0_63674 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[15]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_samples_per_point[15]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73730);
    
    \General_Controller_0/status_bits_1[35]\ : DFN1E1
      port map(D => Pressure_Signal_Debounce_0_low_pressure, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74266, Q => 
        \Data_Hub_Packets_0_status_packet[2]\);
    
    HIEFFPLA_INST_0_58940 : NOR3A
      port map(A => Communications_0_ext_tx_rdy, B => 
        HIEFFPLA_NET_0_74653, C => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74654);
    
    HIEFFPLA_INST_0_56873 : MX2
      port map(A => HIEFFPLA_NET_0_75002, B => 
        HIEFFPLA_NET_0_74930, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75201);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[10]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[10]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[10]\);
    
    HIEFFPLA_INST_0_70805 : AO1A
      port map(A => HIEFFPLA_NET_0_72540, B => 
        HIEFFPLA_NET_0_72009, C => HIEFFPLA_NET_0_72449, Y => 
        HIEFFPLA_NET_0_72461);
    
    HIEFFPLA_INST_0_61320 : NOR2A
      port map(A => HIEFFPLA_NET_0_74210, B => 
        HIEFFPLA_NET_0_74217, Y => HIEFFPLA_NET_0_74218);
    
    \General_Controller_0/sweep_table_write_value[12]\ : DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[12]_net_1\);
    
    HIEFFPLA_INST_0_58112 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_74849);
    
    HIEFFPLA_INST_0_64538 : AND2B
      port map(A => \General_Controller_0/uc_tx_state[12]_net_1\, 
        B => \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73605);
    
    HIEFFPLA_INST_0_60017 : MX2
      port map(A => \Science_0_chan3_data[8]\, B => 
        \Science_0_chan2_data[0]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74473);
    
    \UC_PWR_EN_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => UC_PWR_EN_c, E => \VCC\, DOUT => 
        \UC_PWR_EN_pad/U0/NET1\, EOUT => \UC_PWR_EN_pad/U0/NET2\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[23]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[23]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[23]\);
    
    \Timing_0/s_count[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72056, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_count[0]_net_1\);
    
    HIEFFPLA_INST_0_68701 : OA1C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[0]_net_1\, B
         => HIEFFPLA_NET_0_72668, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_72583);
    
    HIEFFPLA_INST_0_65480 : NOR2A
      port map(A => HIEFFPLA_NET_0_73276, B => 
        \Science_0/ADC_READ_0/cnt2up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73366);
    
    HIEFFPLA_INST_0_71063 : OA1A
      port map(A => HIEFFPLA_NET_0_74284, B => 
        HIEFFPLA_NET_0_74281, C => 
        \General_Controller_0/flight_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74288);
    
    HIEFFPLA_INST_0_62898 : AO1B
      port map(A => HIEFFPLA_NET_0_73918, B => 
        HIEFFPLA_NET_0_73778, C => HIEFFPLA_NET_0_73871, Y => 
        HIEFFPLA_NET_0_73872);
    
    HIEFFPLA_INST_0_63918 : MX2
      port map(A => HIEFFPLA_NET_0_73667, B => 
        HIEFFPLA_NET_0_73660, S => HIEFFPLA_NET_0_73594, Y => 
        HIEFFPLA_NET_0_73690);
    
    HIEFFPLA_INST_0_67840 : AO16
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72790);
    
    HIEFFPLA_INST_0_61210 : OR3A
      port map(A => HIEFFPLA_NET_0_74253, B => 
        \General_Controller_0/state_seconds[3]_net_1\, C => 
        HIEFFPLA_NET_0_74259, Y => HIEFFPLA_NET_0_74249);
    
    HIEFFPLA_INST_0_57873 : AO1
      port map(A => \Science_0_exp_packet_0[78]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75137, Y => HIEFFPLA_NET_0_74919);
    
    HIEFFPLA_INST_0_58058 : AO1
      port map(A => \Sensors_0_gyro_y[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75160, Y => HIEFFPLA_NET_0_74867);
    
    \Science_0/ADC_READ_0/exp_packet_1[77]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[21]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[77]\);
    
    HIEFFPLA_INST_0_65728 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt[0]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73297);
    
    HIEFFPLA_INST_0_69725 : NOR2A
      port map(A => HIEFFPLA_NET_0_72380, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72321);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[21]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[21]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[21]\);
    
    \Communications_0/UART_1/tx_clk_count[7]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75403, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_clk_count_i_0[7]\);
    
    HIEFFPLA_INST_0_66301 : AND2
      port map(A => \Science_0/SWEEP_SPIDER2_0/latch_i_0\, B => 
        \s_clks_net_0[9]\, Y => HIEFFPLA_NET_0_73151);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_11\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[5]\\\\\, CLK => 
        CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_11_Q\);
    
    HIEFFPLA_INST_0_69553 : NOR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        B => HIEFFPLA_NET_0_72375, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72366);
    
    \Science_0/ADC_READ_0/data_a[9]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[9]_net_1\);
    
    HIEFFPLA_INST_0_58450 : NAND2
      port map(A => \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, 
        B => General_Controller_0_en_data_saving, Y => 
        HIEFFPLA_NET_0_74763);
    
    HIEFFPLA_INST_0_56086 : NAND3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[2]\\\\\, B
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[1]\\\\\, 
        C => HIEFFPLA_NET_0_75369, Y => HIEFFPLA_NET_0_75350);
    
    HIEFFPLA_INST_0_68169 : OR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, B
         => CLKINT_1_Y, Y => HIEFFPLA_NET_0_72717);
    
    HIEFFPLA_INST_0_70703 : AND2A
      port map(A => HIEFFPLA_NET_0_72036, B => \s_time[5]\, Y => 
        HIEFFPLA_NET_0_72037);
    
    HIEFFPLA_INST_0_66927 : OA1C
      port map(A => HIEFFPLA_NET_0_72736, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        C => HIEFFPLA_NET_0_72999, Y => HIEFFPLA_NET_0_73003);
    
    HIEFFPLA_INST_0_55561 : NOR3B
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\, B => 
        HIEFFPLA_NET_0_75468, C => 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\, Y => 
        HIEFFPLA_NET_0_75480);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[2]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72217, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[2]_net_1\);
    
    HIEFFPLA_INST_0_69751 : OR3A
      port map(A => HIEFFPLA_NET_0_72314, B => CLKINT_1_Y, C => 
        HIEFFPLA_NET_0_72315, Y => HIEFFPLA_NET_0_72316);
    
    \Science_0/DAC_SET_0/state[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73211, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/state[2]_net_1\);
    
    HIEFFPLA_INST_0_67725 : AND3
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/isSetup_net_1\, 
        C => General_Controller_0_en_sensors, Y => 
        HIEFFPLA_NET_0_72815);
    
    HIEFFPLA_INST_0_66031 : NOR2A
      port map(A => \Science_0/ADC_RESET_0/state[0]_net_1\, B => 
        \Science_0/ADC_RESET_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73232);
    
    HIEFFPLA_INST_0_63188 : AOI1C
      port map(A => HIEFFPLA_NET_0_73913, B => 
        HIEFFPLA_NET_0_73985, C => HIEFFPLA_NET_0_73788, Y => 
        HIEFFPLA_NET_0_73813);
    
    \General_Controller_0/constant_bias_voltage_1[5]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[5]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[5]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[8]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72803, Q => 
        \Sensors_0_mag_x[8]\);
    
    HIEFFPLA_INST_0_58334 : AO1
      port map(A => \Sensors_0_mag_x[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75095, Y => HIEFFPLA_NET_0_74799);
    
    \Timing_0/s_count[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72053, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_count[4]_net_1\);
    
    HIEFFPLA_INST_0_68911 : NOR3B
      port map(A => HIEFFPLA_NET_0_72515, B => 
        HIEFFPLA_NET_0_72486, C => HIEFFPLA_NET_0_72487, Y => 
        HIEFFPLA_NET_0_72524);
    
    HIEFFPLA_INST_0_59079 : NOR3B
      port map(A => HIEFFPLA_NET_0_74448, B => 
        \GS_Readout_0/state[1]_net_1\, C => HIEFFPLA_NET_0_74725, 
        Y => HIEFFPLA_NET_0_74619);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]\ : 
        DFN1P1
      port map(D => HIEFFPLA_NET_0_72210, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\);
    
    HIEFFPLA_INST_0_65126 : AOI1C
      port map(A => HIEFFPLA_NET_0_73465, B => 
        HIEFFPLA_NET_0_73461, C => HIEFFPLA_NET_0_73427, Y => 
        HIEFFPLA_NET_0_73464);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[1]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[1]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[1]\);
    
    HIEFFPLA_INST_0_66455 : NAND3
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        C => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73116);
    
    HIEFFPLA_INST_0_67111 : MX2
      port map(A => HIEFFPLA_NET_0_72917, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[1]\, 
        S => HIEFFPLA_NET_0_72932, Y => HIEFFPLA_NET_0_72962);
    
    HIEFFPLA_INST_0_55764 : AOI1
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\, B => 
        \Communications_0/UART_1/rx_state[0]_net_1\, C => 
        \Communications_0/UART_1/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75429);
    
    \Pressure_Signal_Debounce_0/ms_cnt[4]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73491, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[4]_net_1\);
    
    HIEFFPLA_INST_0_70035 : AND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[5]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72239);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[9]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[9]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[9]\);
    
    HIEFFPLA_INST_0_60635 : MX2
      port map(A => \Science_0_chan3_data[11]\, B => 
        \Science_0_chan2_data[3]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74383);
    
    \Eject_Signal_Debounce_0/state[1]\ : DFN1E1P1
      port map(D => HIEFFPLA_NET_0_74734, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, E => HIEFFPLA_NET_0_72220, Q => 
        \Eject_Signal_Debounce_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_67640 : NOR3B
      port map(A => HIEFFPLA_NET_0_72743, B => 
        HIEFFPLA_NET_0_72885, C => HIEFFPLA_NET_0_72792, Y => 
        HIEFFPLA_NET_0_72835);
    
    HIEFFPLA_INST_0_64476 : OA1C
      port map(A => HIEFFPLA_NET_0_73618, B => 
        HIEFFPLA_NET_0_74323, C => 
        \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73619);
    
    HIEFFPLA_INST_0_64769 : OR3A
      port map(A => HIEFFPLA_NET_0_73542, B => 
        HIEFFPLA_NET_0_73540, C => HIEFFPLA_NET_0_73544, Y => 
        HIEFFPLA_NET_0_73545);
    
    HIEFFPLA_INST_0_58262 : AO1
      port map(A => \Sensors_0_gyro_time[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75109, Y => HIEFFPLA_NET_0_74817);
    
    HIEFFPLA_INST_0_60394 : NOR2A
      port map(A => HIEFFPLA_NET_0_74363, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74421);
    
    HIEFFPLA_INST_0_56124 : AO1
      port map(A => HIEFFPLA_NET_0_75361, B => 
        HIEFFPLA_NET_0_75311, C => HIEFFPLA_NET_0_75340, Y => 
        HIEFFPLA_NET_0_75341);
    
    \Data_Saving_0/Packet_Saver_0/data_out[22]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75222, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[22]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[17]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72280, Q => \Sensors_0_pressure_raw[17]\);
    
    \General_Controller_0/old_1Hz\ : DFN1P1
      port map(D => \AFLSDF_INV_25\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => \General_Controller_0/old_1Hz_i_0\);
    
    HIEFFPLA_INST_0_69446 : NOR2A
      port map(A => HIEFFPLA_NET_0_72430, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_i2c_addr[0]\, 
        Y => HIEFFPLA_NET_0_72386);
    
    \Communications_0/UART_1/rx_clk_count[23]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75465, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75443, Q => 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[57]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[1]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[57]\);
    
    HIEFFPLA_INST_0_68853 : AND2B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, B
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72539);
    
    \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_72695, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\);
    
    \FMC_DA_pad[3]/U0/U0\ : IOPAD_TRI
      port map(D => \FMC_DA_pad[3]/U0/NET1\, E => 
        \FMC_DA_pad[3]/U0/NET2\, PAD => FMC_DA(3));
    
    \Communications_0/UART_0/tx_byte[6]\ : DFN1E1
      port map(D => \GS_Readout_0_send[6]\, CLK => CLKINT_0_Y_0, 
        E => HIEFFPLA_NET_0_75504, Q => 
        \Communications_0/UART_0/tx_byte[6]_net_1\);
    
    HIEFFPLA_INST_0_62333 : AO1C
      port map(A => HIEFFPLA_NET_0_73796, B => 
        \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74003);
    
    \General_Controller_0/flight_state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74291, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/flight_state[1]_net_1\);
    
    \General_Controller_0/st_waddr[6]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_waddr[6]\);
    
    HIEFFPLA_INST_0_66724 : NOR3A
      port map(A => HIEFFPLA_NET_0_73053, B => 
        HIEFFPLA_NET_0_73039, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73054);
    
    HIEFFPLA_INST_0_55623 : AND2
      port map(A => HIEFFPLA_NET_0_75470, B => 
        \Communications_0/UART_1/rx_clk_count[26]_net_1\, Y => 
        HIEFFPLA_NET_0_75462);
    
    HIEFFPLA_INST_0_63133 : NAND3C
      port map(A => HIEFFPLA_NET_0_73821, B => 
        HIEFFPLA_NET_0_73839, C => HIEFFPLA_NET_0_73845, Y => 
        HIEFFPLA_NET_0_73822);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/data_out_1[1]\ : 
        DFN1E0C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72270, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[1]\);
    
    \General_Controller_0/state_seconds[17]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74230, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[17]_net_1\);
    
    \General_Controller_0/st_wdata[13]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[13]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[13]\);
    
    HIEFFPLA_INST_0_60179 : AND3
      port map(A => HIEFFPLA_NET_0_74637, B => 
        HIEFFPLA_NET_0_74654, C => HIEFFPLA_NET_0_74441, Y => 
        HIEFFPLA_NET_0_74449);
    
    \Communications_0/UART_0/rx_count[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75561, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/rx_count[0]_net_1\);
    
    HIEFFPLA_INST_0_70732 : AX1C
      port map(A => HIEFFPLA_NET_0_72032, B => 
        HIEFFPLA_NET_0_72029, C => \Timing_0/m_count[7]_net_1\, Y
         => HIEFFPLA_NET_0_72028);
    
    HIEFFPLA_INST_0_69531 : NOR3A
      port map(A => HIEFFPLA_NET_0_72369, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_72345, Y => HIEFFPLA_NET_0_72370);
    
    HIEFFPLA_INST_0_58120 : AO1
      port map(A => \Science_0_exp_packet_0[38]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_75128, Y => HIEFFPLA_NET_0_74846);
    
    \L2WR_pad/U0/U0\ : IOPAD_TRI
      port map(D => \L2WR_pad/U0/NET1\, E => \L2WR_pad/U0/NET2\, 
        PAD => L2WR);
    
    HIEFFPLA_INST_0_60568 : AND2
      port map(A => HIEFFPLA_NET_0_74517, B => 
        HIEFFPLA_NET_0_74459, Y => HIEFFPLA_NET_0_74394);
    
    \Data_Saving_0/Packet_Saver_0/data_out[14]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75231, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[14]\);
    
    HIEFFPLA_INST_0_65640 : NAND2B
      port map(A => \Science_0/ADC_READ_0/cnt4dn[6]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt4dn[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73320);
    
    \General_Controller_0/status_bits_1[36]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74208, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[3]\);
    
    HIEFFPLA_INST_0_56496 : XNOR2
      port map(A => HIEFFPLA_NET_0_75350, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, Y
         => HIEFFPLA_NET_0_75264);
    
    \General_Controller_0/unit_id[2]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73990, Q => 
        \General_Controller_0_unit_id[2]\);
    
    HIEFFPLA_INST_0_58372 : AO1
      port map(A => \Sensors_0_mag_time[15]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75115, Y => HIEFFPLA_NET_0_74789);
    
    \Science_0/ADC_READ_0/chan7_data[8]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[8]\);
    
    HIEFFPLA_INST_0_70746 : AND2
      port map(A => HIEFFPLA_NET_0_72021, B => 
        \Timing_0/s_count[4]_net_1\, Y => HIEFFPLA_NET_0_72024);
    
    HIEFFPLA_INST_0_69280 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, C
         => HIEFFPLA_NET_0_72540, Y => HIEFFPLA_NET_0_72431);
    
    HIEFFPLA_INST_0_62504 : AOI1
      port map(A => HIEFFPLA_NET_0_73864, B => 
        HIEFFPLA_NET_0_73987, C => HIEFFPLA_NET_0_74036, Y => 
        HIEFFPLA_NET_0_73969);
    
    HIEFFPLA_INST_0_68488 : NOR2A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\, B
         => \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_72639);
    
    HIEFFPLA_INST_0_55217 : XNOR2
      port map(A => \Communications_0/UART_0/rx_count[1]_net_1\, 
        B => \Communications_0/UART_0/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75558);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRYSYNC[6]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_16_Q\, 
        CLK => CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[6]\\\\\);
    
    \UC_CONSOLE_EN_pad/U0/U1\ : IOIN_IB
      port map(YIN => \UC_CONSOLE_EN_pad/U0/NET1\, Y => 
        UC_CONSOLE_EN_c);
    
    HIEFFPLA_INST_0_57185 : AND2
      port map(A => \Sensors_0_pressure_time[22]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75136);
    
    HIEFFPLA_INST_0_59098 : AO1A
      port map(A => HIEFFPLA_NET_0_74382, B => 
        \GS_Readout_0/state[1]_net_1\, C => HIEFFPLA_NET_0_74594, 
        Y => HIEFFPLA_NET_0_74613);
    
    HIEFFPLA_INST_0_58427 : OA1C
      port map(A => HIEFFPLA_NET_0_74772, B => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, C => 
        HIEFFPLA_NET_0_74769, Y => HIEFFPLA_NET_0_74770);
    
    HIEFFPLA_INST_0_57214 : AND2
      port map(A => \Sensors_0_acc_time[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, Y
         => HIEFFPLA_NET_0_75127);
    
    HIEFFPLA_INST_0_67938 : MX2
      port map(A => HIEFFPLA_NET_0_72755, B => 
        HIEFFPLA_NET_0_72748, S => HIEFFPLA_NET_0_72878, Y => 
        HIEFFPLA_NET_0_72769);
    
    HIEFFPLA_INST_0_57967 : AO1
      port map(A => \Science_0_exp_packet_0[24]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74788, Y => HIEFFPLA_NET_0_74891);
    
    \GS_Readout_0/state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74612, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/state[1]_net_1\);
    
    \General_Controller_0/sweep_table_sample_skip[8]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[8]_net_1\);
    
    \Science_0/DAC_SET_0/ADR[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73228, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[6]\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72293, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72221, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[6]_net_1\);
    
    HIEFFPLA_INST_0_68683 : NOR3A
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, C
         => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72588);
    
    HIEFFPLA_INST_0_65606 : NOR3B
      port map(A => HIEFFPLA_NET_0_73338, B => 
        \Science_0/ADC_READ_0/cnt3up[2]_net_1\, C => 
        HIEFFPLA_NET_0_73330, Y => HIEFFPLA_NET_0_73332);
    
    HIEFFPLA_INST_0_58677 : AND3C
      port map(A => HIEFFPLA_NET_0_74626, B => 
        HIEFFPLA_NET_0_74648, C => HIEFFPLA_NET_0_74659, Y => 
        HIEFFPLA_NET_0_74706);
    
    HIEFFPLA_INST_0_64185 : AO1A
      port map(A => \General_Controller_0/uc_tx_state[14]_net_1\, 
        B => HIEFFPLA_NET_0_73750, C => 
        \General_Controller_0/uc_tx_state[12]_net_1\, Y => 
        HIEFFPLA_NET_0_73654);
    
    \Timing_0/s_time[5]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72049, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \s_time[5]\);
    
    HIEFFPLA_INST_0_64819 : AND2
      port map(A => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73533);
    
    HIEFFPLA_INST_0_66180 : NOR2A
      port map(A => \Science_0/DAC_SET_0/state[3]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73186);
    
    HIEFFPLA_INST_0_65203 : AX1C
      port map(A => HIEFFPLA_NET_0_73444, B => 
        HIEFFPLA_NET_0_73442, C => 
        \Pressure_Signal_Debounce_0/ms_cnt[8]_net_1\, Y => 
        HIEFFPLA_NET_0_73446);
    
    HIEFFPLA_INST_0_66036 : NAND2B
      port map(A => \Science_0/DAC_SET_0/ADR[0]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73230);
    
    HIEFFPLA_INST_0_60787 : MX2
      port map(A => HIEFFPLA_NET_0_74563, B => 
        HIEFFPLA_NET_0_74554, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74358);
    
    HIEFFPLA_INST_0_56295 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[2]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[1]\\\\\, Y => 
        HIEFFPLA_NET_0_75316);
    
    AFLSDF_INV_20 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_20\);
    
    HIEFFPLA_INST_0_57200 : AO1
      port map(A => \Sensors_0_pressure_time[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75091, Y => HIEFFPLA_NET_0_75132);
    
    \UC_I2C4_SCL_pad/U0/U0\ : IOPAD_IN
      port map(PAD => UC_I2C4_SCL, Y => \UC_I2C4_SCL_pad/U0/NET1\);
    
    HIEFFPLA_INST_0_56806 : MX2
      port map(A => HIEFFPLA_NET_0_75171, B => 
        HIEFFPLA_NET_0_75025, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75208);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/temp[1]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72907, Q => 
        \Sensors_0_acc_temp[1]\);
    
    HIEFFPLA_INST_0_66525 : AO1
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\, 
        B => ACCE_SCL_c, C => HIEFFPLA_NET_0_73048, Y => 
        HIEFFPLA_NET_0_73102);
    
    HIEFFPLA_INST_0_62227 : AND3
      port map(A => HIEFFPLA_NET_0_74113, B => 
        HIEFFPLA_NET_0_74092, C => HIEFFPLA_NET_0_73986, Y => 
        HIEFFPLA_NET_0_74025);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[11]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72800, Q => 
        \Sensors_0_acc_x[11]\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]\ : 
        DFN0E0
      port map(D => HIEFFPLA_NET_0_73105, CLK => 
        ClockDivs_0_clk_800kHz, E => HIEFFPLA_NET_0_73056, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\);
    
    HIEFFPLA_INST_0_69766 : NOR3A
      port map(A => HIEFFPLA_NET_0_72278, B => 
        HIEFFPLA_NET_0_72308, C => HIEFFPLA_NET_0_72305, Y => 
        HIEFFPLA_NET_0_72312);
    
    HIEFFPLA_INST_0_63018 : AND3
      port map(A => HIEFFPLA_NET_0_74077, B => 
        HIEFFPLA_NET_0_74105, C => HIEFFPLA_NET_0_73840, Y => 
        HIEFFPLA_NET_0_73846);
    
    HIEFFPLA_INST_0_59997 : MX2
      port map(A => \Science_0_chan1_data[3]\, B => 
        \Science_0_chan1_data[7]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74476);
    
    HIEFFPLA_INST_0_70499 : XOR2
      port map(A => HIEFFPLA_NET_0_72121, B => 
        \Timekeeper_0_milliseconds[17]\, Y => 
        HIEFFPLA_NET_0_72108);
    
    HIEFFPLA_INST_0_61832 : MX2
      port map(A => HIEFFPLA_NET_0_74082, B => 
        HIEFFPLA_NET_0_74108, S => 
        \General_Controller_0/uc_rx_byte_0[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74119);
    
    \General_Controller_0/uc_tx_state[6]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73567, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[6]_net_1\);
    
    HIEFFPLA_INST_0_64449 : NOR3B
      port map(A => HIEFFPLA_NET_0_74018, B => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, C => 
        HIEFFPLA_NET_0_73897, Y => HIEFFPLA_NET_0_73624);
    
    HIEFFPLA_INST_0_64287 : MX2
      port map(A => HIEFFPLA_NET_0_73729, B => 
        HIEFFPLA_NET_0_73721, S => HIEFFPLA_NET_0_73619, Y => 
        HIEFFPLA_NET_0_73641);
    
    \General_Controller_0/sweep_table_read_value[5]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74159, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[5]_net_1\);
    
    HIEFFPLA_INST_0_60542 : MX2
      port map(A => HIEFFPLA_NET_0_74455, B => 
        HIEFFPLA_NET_0_74488, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74398);
    
    HIEFFPLA_INST_0_58090 : AND2
      port map(A => \ch3_data_net_0[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_74857);
    
    HIEFFPLA_INST_0_58041 : AO1
      port map(A => \Sensors_0_mag_x[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_75143, Y => HIEFFPLA_NET_0_74870);
    
    \Science_0/ADC_READ_0/exp_packet_1[32]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[16]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[32]\);
    
    HIEFFPLA_INST_0_60159 : MX2
      port map(A => \Science_0_chan3_data[3]\, B => 
        \Science_0_chan3_data[7]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74452);
    
    \Timekeeper_0/milliseconds[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72116, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timekeeper_0_milliseconds[0]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[16]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72282, Q => 
        \Sensors_0_pressure_temp_raw[16]\);
    
    HIEFFPLA_INST_0_62107 : AO1
      port map(A => 
        \General_Controller_0/uc_rx_prev_state[1]_net_1\, B => 
        HIEFFPLA_NET_0_73943, C => HIEFFPLA_NET_0_74049, Y => 
        HIEFFPLA_NET_0_74051);
    
    HIEFFPLA_INST_0_61618 : AND2
      port map(A => HIEFFPLA_NET_0_74181, B => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74173);
    
    \Science_0/SET_LP_GAIN_0/state[2]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73157, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/state_i_0[2]\);
    
    \General_Controller_0/state_seconds[9]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74218, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[9]_net_1\);
    
    \General_Controller_0/status_bits_1[58]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74188, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[58]\);
    
    \Science_0/SET_LP_GAIN_0/L3WR\ : DFN0C1
      port map(D => \Science_0/SET_LP_GAIN_0/state_i_0[1]\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => L3WR_c);
    
    HIEFFPLA_INST_0_58423 : AND3C
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\, B => 
        \Data_Saving_0/Packet_Saver_0/acc_flag_net_1\, C => 
        \Data_Saving_0/Packet_Saver_0/mag_flag_net_1\, Y => 
        HIEFFPLA_NET_0_74771);
    
    HIEFFPLA_INST_0_56436 : MX2
      port map(A => \FMC_DA_c[5]\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[5]\\\\\, S => 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\, Y => 
        HIEFFPLA_NET_0_75282);
    
    \General_Controller_0/gs_id[1]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73922, Q => 
        \General_Controller_0_gs_id[1]\);
    
    HIEFFPLA_INST_0_64806 : AX1C
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        HIEFFPLA_NET_0_74013, C => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73537);
    
    HIEFFPLA_INST_0_70052 : NOR2A
      port map(A => HIEFFPLA_NET_0_72233, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        Y => HIEFFPLA_NET_0_72234);
    
    HIEFFPLA_INST_0_70090 : NAND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]_net_1\, 
        B => \Sensors_0/Pressure_Sensor_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72223);
    
    HIEFFPLA_INST_0_62641 : AND3B
      port map(A => HIEFFPLA_NET_0_73811, B => 
        HIEFFPLA_NET_0_73889, C => HIEFFPLA_NET_0_73907, Y => 
        HIEFFPLA_NET_0_73939);
    
    HIEFFPLA_INST_0_69893 : AND3
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[2]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72276);
    
    HIEFFPLA_INST_0_60063 : MX2
      port map(A => \Science_0_chan0_data[5]\, B => 
        \Science_0_chan0_data[9]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74467);
    
    HIEFFPLA_INST_0_69718 : AOI1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        C => HIEFFPLA_NET_0_72410, Y => HIEFFPLA_NET_0_72322);
    
    HIEFFPLA_INST_0_58729 : AND3
      port map(A => HIEFFPLA_NET_0_74692, B => 
        HIEFFPLA_NET_0_74459, C => HIEFFPLA_NET_0_74496, Y => 
        HIEFFPLA_NET_0_74696);
    
    HIEFFPLA_INST_0_64604 : AO1A
      port map(A => 
        \General_Controller_0/uc_tx_substate[2]_net_1\, B => 
        HIEFFPLA_NET_0_73589, C => HIEFFPLA_NET_0_73554, Y => 
        HIEFFPLA_NET_0_73590);
    
    HIEFFPLA_INST_0_58326 : AO1
      port map(A => \Sensors_0_mag_x[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75083, Y => HIEFFPLA_NET_0_74801);
    
    HIEFFPLA_INST_0_57853 : AO1
      port map(A => \Science_0_exp_packet_0[76]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75139, Y => HIEFFPLA_NET_0_74925);
    
    \ACST_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => \VCC\, E => \VCC\, DOUT => \ACST_pad/U0/NET1\, 
        EOUT => \ACST_pad/U0/NET2\);
    
    \Science_0/ADC_READ_0/data_a[4]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[3]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[4]_net_1\);
    
    HIEFFPLA_INST_0_66242 : MX2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G3[0]_net_1\, B
         => \Science_0/ADC_READ_0_G3[0]\, S => 
        \Science_0/SET_LP_GAIN_0/state[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73169);
    
    HIEFFPLA_INST_0_62979 : NAND3C
      port map(A => HIEFFPLA_NET_0_73852, B => 
        HIEFFPLA_NET_0_73844, C => HIEFFPLA_NET_0_73836, Y => 
        HIEFFPLA_NET_0_73853);
    
    \Science_0/ADC_READ_0/data_a[15]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[15]_net_1\);
    
    HIEFFPLA_INST_0_55515 : NOR3B
      port map(A => HIEFFPLA_NET_0_75483, B => 
        HIEFFPLA_NET_0_75488, C => 
        \Communications_0/UART_1/rx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75491);
    
    HIEFFPLA_INST_0_68814 : AND3
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, B
         => HIEFFPLA_NET_0_72487, C => 
        \Sensors_0/Gyro_0/I2C_Master_0_write_done\, Y => 
        HIEFFPLA_NET_0_72550);
    
    \General_Controller_0/state_seconds[16]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74232, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[16]_net_1\);
    
    \General_Controller_0/sweep_table_step_id[2]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73926, Q => 
        \General_Controller_0/sweep_table_step_id[2]_net_1\);
    
    \General_Controller_0/constant_bias_voltage_1[4]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[4]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[4]_net_1\);
    
    HIEFFPLA_INST_0_68625 : NOR3A
      port map(A => HIEFFPLA_NET_0_72592, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, C
         => \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72603);
    
    HIEFFPLA_INST_0_56019 : XA1A
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[8]\\\\\, B => 
        HIEFFPLA_NET_0_75267, C => HIEFFPLA_NET_0_75356, Y => 
        HIEFFPLA_NET_0_75368);
    
    HIEFFPLA_INST_0_71013 : OA1C
      port map(A => \I2C_PassThrough_0/state[0]_net_1\, B => 
        HIEFFPLA_NET_0_73518, C => \I2C_PassThrough_0.state[3]\, 
        Y => HIEFFPLA_NET_0_71989);
    
    HIEFFPLA_INST_0_69509 : NOR3B
      port map(A => HIEFFPLA_NET_0_72372, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72374);
    
    HIEFFPLA_INST_0_68339 : NAND3A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, C => 
        GYRO_SCL_c, Y => HIEFFPLA_NET_0_72678);
    
    HIEFFPLA_INST_0_58686 : NAND3B
      port map(A => HIEFFPLA_NET_0_74648, B => 
        HIEFFPLA_NET_0_74659, C => HIEFFPLA_NET_0_74668, Y => 
        HIEFFPLA_NET_0_74704);
    
    HIEFFPLA_INST_0_65836 : MX2
      port map(A => HIEFFPLA_NET_0_73270, B => 
        HIEFFPLA_NET_0_73268, S => 
        \Science_0/ADC_READ_0/chan[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73272);
    
    HIEFFPLA_INST_0_65285 : OR3A
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, B => 
        \Science_0/ADC_READ_0/chan[0]_net_1\, C => 
        HIEFFPLA_NET_0_73243, Y => HIEFFPLA_NET_0_73423);
    
    HIEFFPLA_INST_0_55391 : XO1A
      port map(A => HIEFFPLA_NET_0_75536, B => 
        \Communications_0/UART_0/tx_clk_count_i_0[3]\, C => 
        HIEFFPLA_NET_0_75527, Y => HIEFFPLA_NET_0_75523);
    
    \General_Controller_0/sweep_table_points[1]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[1]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[1]_net_1\);
    
    HIEFFPLA_INST_0_60426 : MX2
      port map(A => \Sensors_0_acc_z[7]\, B => 
        \Sensors_0_acc_z[11]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74417);
    
    HIEFFPLA_INST_0_61140 : AND3A
      port map(A => CLKINT_1_Y, B => \s_clks_net_0[18]\, C => 
        \General_Controller_0/old_status_packet_clk_i_0\, Y => 
        HIEFFPLA_NET_0_74266);
    
    \General_Controller_0/temp_first_byte[2]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73872, Q => 
        \General_Controller_0/temp_first_byte[2]_net_1\);
    
    HIEFFPLA_INST_0_68827 : AO1A
      port map(A => HIEFFPLA_NET_0_72540, B => 
        HIEFFPLA_NET_0_72542, C => HIEFFPLA_NET_0_72476, Y => 
        HIEFFPLA_NET_0_72547);
    
    HIEFFPLA_INST_0_56367 : XNOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, B
         => HIEFFPLA_NET_0_75370, Y => HIEFFPLA_NET_0_75299);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_1\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_72378, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72348, Q => 
        \Sensors_0.Pressure_Sensor_0.I2C_Master_0.sda_1\);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]\ : 
        DFN0E1
      port map(D => HIEFFPLA_NET_0_72387, CLK => 
        ClockDivs_0_clk_800kHz, E => HIEFFPLA_NET_0_72354, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[1]_net_1\);
    
    HIEFFPLA_INST_0_67420 : AND3
      port map(A => HIEFFPLA_NET_0_72935, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72886);
    
    HIEFFPLA_INST_0_67093 : NOR2A
      port map(A => HIEFFPLA_NET_0_72961, B => 
        HIEFFPLA_NET_0_72964, Y => HIEFFPLA_NET_0_72965);
    
    HIEFFPLA_INST_0_58385 : AO1
      port map(A => \Sensors_0_gyro_x[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74782, Y => HIEFFPLA_NET_0_74783);
    
    HIEFFPLA_INST_0_55758 : NOR3A
      port map(A => HIEFFPLA_NET_0_75468, B => 
        \Communications_0/UART_1/rx_state[1]_net_1\, C => 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\, Y => 
        HIEFFPLA_NET_0_75431);
    
    \I2C_PassThrough_0/state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73512, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \I2C_PassThrough_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_63927 : AO1
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[14]_net_1\, 
        B => HIEFFPLA_NET_0_73579, C => HIEFFPLA_NET_0_73688, Y
         => HIEFFPLA_NET_0_73689);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[14]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72281, Q => \Sensors_0_pressure_raw[14]\);
    
    HIEFFPLA_INST_0_55697 : NOR2A
      port map(A => General_Controller_0_uc_oen, B => 
        \Communications_0/UART_1/rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75445);
    
    HIEFFPLA_INST_0_65956 : NAND3
      port map(A => \Science_0/ADC_READ_0_G3[0]\, B => 
        \Science_0/ADC_READ_0/cnt3up[4]_net_1\, C => 
        HIEFFPLA_NET_0_73276, Y => HIEFFPLA_NET_0_73252);
    
    HIEFFPLA_INST_0_55607 : NAND2B
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[29]_net_1\, B => 
        \Communications_0/UART_1/rx_clk_count[28]_net_1\, Y => 
        HIEFFPLA_NET_0_75466);
    
    HIEFFPLA_INST_0_61785 : AX1C
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[3]_net_1\, B
         => HIEFFPLA_NET_0_74148, C => 
        \General_Controller_0/sweep_table_sweep_cnt[4]_net_1\, Y
         => HIEFFPLA_NET_0_74134);
    
    \Communications_0/UART_0/rx_clk_count[30]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75569, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75554, Q => 
        \Communications_0/UART_0/rx_clk_count[30]_net_1\);
    
    \Communications_0/UART_1/tx_clk_count[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75410, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_clk_count[1]_net_1\);
    
    HIEFFPLA_INST_0_65395 : XOR2
      port map(A => \Science_0/ADC_READ_0/cnt1up[3]_net_1\, B => 
        HIEFFPLA_NET_0_73388, Y => HIEFFPLA_NET_0_73390);
    
    HIEFFPLA_INST_0_57290 : AND2
      port map(A => \Sensors_0_gyro_time[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75090);
    
    HIEFFPLA_INST_0_65305 : NAND2B
      port map(A => \Science_0/ADC_READ_0/cnt1dn[2]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt1dn[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73416);
    
    HIEFFPLA_INST_0_56300 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, B
         => HIEFFPLA_NET_0_75370, C => HIEFFPLA_NET_0_75312, Y
         => HIEFFPLA_NET_0_75314);
    
    HIEFFPLA_INST_0_62187 : AOI1D
      port map(A => \General_Controller_0/uc_rx_state_0[1]_net_1\, 
        B => HIEFFPLA_NET_0_73888, C => HIEFFPLA_NET_0_73785, Y
         => HIEFFPLA_NET_0_74034);
    
    HIEFFPLA_INST_0_69072 : AO1
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        B => \Sensors_0/Gyro_0/state[8]\, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        Y => HIEFFPLA_NET_0_72477);
    
    \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[2]\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72686, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72618, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[2]_net_1\);
    
    HIEFFPLA_INST_0_56847 : MX2
      port map(A => HIEFFPLA_NET_0_75166, B => 
        HIEFFPLA_NET_0_75013, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75204);
    
    HIEFFPLA_INST_0_57157 : AND2
      port map(A => \Sensors_0_pressure_time[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, Y
         => HIEFFPLA_NET_0_75148);
    
    \Communications_0/UART_0/recv[5]\ : DFN1E1C1
      port map(D => \Communications_0/UART_0/rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75551, Q => 
        \Communications_0/UART_0_recv[5]\);
    
    HIEFFPLA_INST_0_70142 : AND3C
      port map(A => HIEFFPLA_NET_0_72204, B => 
        HIEFFPLA_NET_0_72190, C => HIEFFPLA_NET_0_72182, Y => 
        HIEFFPLA_NET_0_72210);
    
    \General_Controller_0/sweep_table_read_value[7]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74157, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[7]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[2]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[2]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[2]\);
    
    \Science_0/ADC_READ_0/cnt2dn[5]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73371, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2dn[5]_net_1\);
    
    HIEFFPLA_INST_0_70431 : AX1C
      port map(A => \Timekeeper_0_microseconds[3]\, B => 
        HIEFFPLA_NET_0_72154, C => \Timekeeper_0_microseconds[4]\, 
        Y => HIEFFPLA_NET_0_72133);
    
    HIEFFPLA_INST_0_61328 : NOR2A
      port map(A => 
        \General_Controller_0/state_seconds[10]_net_1\, B => 
        HIEFFPLA_NET_0_74241, Y => HIEFFPLA_NET_0_74216);
    
    HIEFFPLA_INST_0_70720 : AND3
      port map(A => \Timing_0/m_count[0]_net_1\, B => 
        \Timing_0/m_count[1]_net_1\, C => 
        \Timing_0/m_count[2]_net_1\, Y => HIEFFPLA_NET_0_72032);
    
    HIEFFPLA_INST_0_70525 : AX1C
      port map(A => \Timekeeper_0_milliseconds[5]\, B => 
        HIEFFPLA_NET_0_72117, C => \Timekeeper_0_milliseconds[6]\, 
        Y => HIEFFPLA_NET_0_72096);
    
    \Timing_0/m_time[5]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72062, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_time[5]_net_1\);
    
    HIEFFPLA_INST_0_56283 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[2]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[1]\\\\\, C => 
        HIEFFPLA_NET_0_75323, Y => HIEFFPLA_NET_0_75319);
    
    \General_Controller_0/st_raddr[5]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[5]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73979, Q => 
        \General_Controller_0_st_raddr_1[5]\);
    
    HIEFFPLA_INST_0_63249 : AO1
      port map(A => HIEFFPLA_NET_0_73951, B => 
        HIEFFPLA_NET_0_73901, C => HIEFFPLA_NET_0_73798, Y => 
        HIEFFPLA_NET_0_73799);
    
    HIEFFPLA_INST_0_59048 : OA1A
      port map(A => HIEFFPLA_NET_0_74490, B => 
        HIEFFPLA_NET_0_74725, C => \GS_Readout_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_74627);
    
    \Pressure_Signal_Debounce_0/ms_cnt[8]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73485, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[8]_net_1\);
    
    HIEFFPLA_INST_0_63710 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[5]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_nof_steps[5]_net_1\, S
         => \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73724);
    
    \Timekeeper_0/microseconds[19]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72141, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[19]\);
    
    \Science_0/SWEEP_SPIDER2_0/latch\ : DFN1P1
      port map(D => \AFLSDF_INV_26\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => \Science_0/SWEEP_SPIDER2_0/latch_i_0\);
    
    HIEFFPLA_INST_0_69332 : XA1B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\, 
        B => HIEFFPLA_NET_0_72320, C => HIEFFPLA_NET_0_72415, Y
         => HIEFFPLA_NET_0_72416);
    
    HIEFFPLA_INST_0_61240 : XA1C
      port map(A => HIEFFPLA_NET_0_74241, B => 
        \General_Controller_0/state_seconds[10]_net_1\, C => 
        HIEFFPLA_NET_0_74217, Y => HIEFFPLA_NET_0_74239);
    
    HIEFFPLA_INST_0_66074 : AX1
      port map(A => HIEFFPLA_NET_0_73223, B => 
        HIEFFPLA_NET_0_73213, C => 
        \Science_0/DAC_SET_0/cnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73217);
    
    HIEFFPLA_INST_0_61901 : NOR3A
      port map(A => \General_Controller_0/uc_rx_byte[0]_net_1\, B
         => HIEFFPLA_NET_0_74082, C => 
        \General_Controller_0/uc_rx_byte[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74103);
    
    HIEFFPLA_INST_0_62888 : AND3C
      port map(A => HIEFFPLA_NET_0_73873, B => 
        \General_Controller_0/uc_rx_state[0]_net_1\, C => 
        HIEFFPLA_NET_0_73811, Y => HIEFFPLA_NET_0_73874);
    
    HIEFFPLA_INST_0_59515 : MX2
      port map(A => HIEFFPLA_NET_0_74497, B => 
        HIEFFPLA_NET_0_74361, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74543);
    
    \Data_Saving_0/Packet_Saver_0/data_out[29]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75214, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[29]\);
    
    HIEFFPLA_INST_0_69909 : NAND3C
      port map(A => HIEFFPLA_NET_0_72285, B => 
        HIEFFPLA_NET_0_72278, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72269);
    
    CLKINT_2 : CLKINT
      port map(A => FMC_CLK_c, Y => CLKINT_2_Y);
    
    HIEFFPLA_INST_0_57753 : AO1B
      port map(A => \Sensors_0_acc_x[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74952, Y => HIEFFPLA_NET_0_74953);
    
    HIEFFPLA_INST_0_67579 : NOR3B
      port map(A => HIEFFPLA_NET_0_72819, B => 
        HIEFFPLA_NET_0_72817, C => HIEFFPLA_NET_0_72945, Y => 
        HIEFFPLA_NET_0_72848);
    
    HIEFFPLA_INST_0_61892 : AND2
      port map(A => \General_Controller_0/uc_rx_byte[1]_net_1\, B
         => \General_Controller_0/uc_rx_byte[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74107);
    
    HIEFFPLA_INST_0_56995 : NOR3A
      port map(A => HIEFFPLA_NET_0_74960, B => 
        HIEFFPLA_NET_0_75127, C => HIEFFPLA_NET_0_74844, Y => 
        HIEFFPLA_NET_0_75185);
    
    HIEFFPLA_INST_0_65642 : AND3
      port map(A => HIEFFPLA_NET_0_73321, B => 
        HIEFFPLA_NET_0_73325, C => HIEFFPLA_NET_0_73277, Y => 
        HIEFFPLA_NET_0_73319);
    
    HIEFFPLA_INST_0_62447 : NOR3B
      port map(A => HIEFFPLA_NET_0_74037, B => 
        HIEFFPLA_NET_0_73887, C => HIEFFPLA_NET_0_73776, Y => 
        HIEFFPLA_NET_0_73980);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[0]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72276, Q => \Sensors_0_pressure_raw[0]\);
    
    HIEFFPLA_INST_0_58287 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[54]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_74811);
    
    \Data_Saving_0/Packet_Saver_0/ch_0_flag\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_75238, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => 
        General_Controller_0_en_data_saving, Q => 
        \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\);
    
    HIEFFPLA_INST_0_65933 : NAND2B
      port map(A => HIEFFPLA_NET_0_73255, B => 
        HIEFFPLA_NET_0_73256, Y => HIEFFPLA_NET_0_73257);
    
    HIEFFPLA_INST_0_59753 : MX2
      port map(A => HIEFFPLA_NET_0_74532, B => 
        HIEFFPLA_NET_0_74524, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74513);
    
    HIEFFPLA_INST_0_67950 : NOR3B
      port map(A => HIEFFPLA_NET_0_72889, B => 
        HIEFFPLA_NET_0_72790, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72768);
    
    HIEFFPLA_INST_0_62815 : OR3B
      port map(A => HIEFFPLA_NET_0_73903, B => 
        HIEFFPLA_NET_0_73894, C => HIEFFPLA_NET_0_73795, Y => 
        HIEFFPLA_NET_0_73895);
    
    HIEFFPLA_INST_0_57100 : MX2
      port map(A => HIEFFPLA_NET_0_74936, B => 
        HIEFFPLA_NET_0_74881, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75167);
    
    \Communications_0/UART_0/rx_byte[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75380, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75606, Q => 
        \Communications_0/UART_0/rx_byte[6]_net_1\);
    
    \Timekeeper_0/milliseconds[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72100, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[2]\);
    
    HIEFFPLA_INST_0_69950 : AO1A
      port map(A => HIEFFPLA_NET_0_72250, B => 
        HIEFFPLA_NET_0_72248, C => HIEFFPLA_NET_0_72255, Y => 
        HIEFFPLA_NET_0_72261);
    
    HIEFFPLA_INST_0_59947 : NOR3A
      port map(A => HIEFFPLA_NET_0_74408, B => 
        HIEFFPLA_NET_0_74360, C => HIEFFPLA_NET_0_74634, Y => 
        HIEFFPLA_NET_0_74484);
    
    \General_Controller_0/sweep_table_sample_skip[0]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[0]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[0]_net_1\);
    
    HIEFFPLA_INST_0_67404 : OR3A
      port map(A => HIEFFPLA_NET_0_72799, B => 
        HIEFFPLA_NET_0_72877, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72890);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[13]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72553, Q => 
        \Sensors_0_gyro_x[13]\);
    
    HIEFFPLA_INST_0_68787 : AO1A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, B
         => HIEFFPLA_NET_0_72539, C => HIEFFPLA_NET_0_72561, Y
         => HIEFFPLA_NET_0_72562);
    
    HIEFFPLA_INST_0_64899 : AOI1C
      port map(A => \I2C_PassThrough_0/state[1]_net_1\, B => 
        \I2C_PassThrough_0/state[0]_net_1\, C => CLKINT_1_Y, Y
         => HIEFFPLA_NET_0_73514);
    
    HIEFFPLA_INST_0_61633 : MX2
      port map(A => \SweepTable_0_RD[10]\, B => 
        \SweepTable_1_RD[10]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74169);
    
    \PRESSURE_SCL_pad/U0/U0\ : IOPAD_TRI
      port map(D => \PRESSURE_SCL_pad/U0/NET1\, E => 
        \PRESSURE_SCL_pad/U0/NET2\, PAD => PRESSURE_SCL);
    
    HIEFFPLA_INST_0_59460 : MX2
      port map(A => HIEFFPLA_NET_0_74418, B => 
        HIEFFPLA_NET_0_74437, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74551);
    
    HIEFFPLA_INST_0_56248 : XOR3
      port map(A => HIEFFPLA_NET_0_75322, B => 
        HIEFFPLA_NET_0_75319, C => HIEFFPLA_NET_0_75264, Y => 
        HIEFFPLA_NET_0_75325);
    
    HIEFFPLA_INST_0_65121 : NAND3
      port map(A => \Sensors_0_pressure_raw[10]\, B => 
        \Sensors_0_pressure_raw[13]\, C => 
        \Sensors_0_pressure_raw[12]\, Y => HIEFFPLA_NET_0_73466);
    
    \Data_Saving_0/Packet_Saver_0/word_cnt[0]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_74762, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[43]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[9]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[43]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/num_bytes_1[0]\ : 
        DFN1E0C1
      port map(D => HIEFFPLA_NET_0_72291, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72232, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_num_bytes[0]\);
    
    HIEFFPLA_INST_0_62172 : AND3A
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74037);
    
    HIEFFPLA_INST_0_70602 : AND3
      port map(A => \Timing_0/m_time[4]_net_1\, B => 
        \Timing_0/m_time[5]_net_1\, C => HIEFFPLA_NET_0_72070, Y
         => HIEFFPLA_NET_0_72068);
    
    HIEFFPLA_INST_0_65931 : AO1B
      port map(A => HIEFFPLA_NET_0_73276, B => 
        \Science_0/ADC_READ_0/cnt2up[4]_net_1\, C => 
        \Science_0/ADC_READ_0_G2[0]\, Y => HIEFFPLA_NET_0_73258);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[0]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[0]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[0]\);
    
    \Timing_0/s_count[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72054, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_count[3]_net_1\);
    
    HIEFFPLA_INST_0_55761 : AND2B
      port map(A => HIEFFPLA_NET_0_75482, B => 
        \Communications_0/UART_1/rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75430);
    
    \Science_0/ADC_READ_0/chan3_data[7]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[7]\);
    
    HIEFFPLA_INST_0_67276 : NOR3B
      port map(A => HIEFFPLA_NET_0_72760, B => 
        HIEFFPLA_NET_0_72882, C => HIEFFPLA_NET_0_72717, Y => 
        HIEFFPLA_NET_0_72920);
    
    \General_Controller_0/sweep_table_samples_per_point[12]\ : 
        DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[12]_net_1\);
    
    HIEFFPLA_INST_0_70484 : AX1
      port map(A => \Timekeeper_0/old_1kHz_net_1\, B => 
        \m_time[7]\, C => \Timekeeper_0_milliseconds[0]\, Y => 
        HIEFFPLA_NET_0_72116);
    
    HIEFFPLA_INST_0_70567 : XA1B
      port map(A => HIEFFPLA_NET_0_72032, B => 
        \Timing_0/m_count[3]_net_1\, C => HIEFFPLA_NET_0_72083, Y
         => HIEFFPLA_NET_0_72077);
    
    HIEFFPLA_INST_0_59090 : NOR3B
      port map(A => HIEFFPLA_NET_0_74443, B => 
        \GS_Readout_0/state[4]_net_1\, C => HIEFFPLA_NET_0_74725, 
        Y => HIEFFPLA_NET_0_74615);
    
    \Science_0/ADC_READ_0/data_b[14]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[14]_net_1\);
    
    \Science_0/SET_LP_GAIN_0/state[0]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73161, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/state_i_0[0]\);
    
    HIEFFPLA_INST_0_67979 : NAND3B
      port map(A => HIEFFPLA_NET_0_72935, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_72881, Y => HIEFFPLA_NET_0_72763);
    
    HIEFFPLA_INST_0_59772 : MX2
      port map(A => \Science_0_chan1_data[1]\, B => 
        \Science_0_chan1_data[5]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74511);
    
    HIEFFPLA_INST_0_70048 : OR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        B => HIEFFPLA_NET_0_72242, C => HIEFFPLA_NET_0_72229, Y
         => HIEFFPLA_NET_0_72235);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[22]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72280, Q => \Sensors_0_pressure_raw[22]\);
    
    HIEFFPLA_INST_0_64637 : AND3B
      port map(A => \General_Controller_0/uc_tx_state[15]_net_1\, 
        B => \General_Controller_0/uc_tx_state[14]_net_1\, C => 
        HIEFFPLA_NET_0_73605, Y => HIEFFPLA_NET_0_73580);
    
    \Science_0/ADC_READ_0/chan4_data[3]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[3]\);
    
    HIEFFPLA_INST_0_63110 : NOR3B
      port map(A => HIEFFPLA_NET_0_74091, B => 
        HIEFFPLA_NET_0_73841, C => HIEFFPLA_NET_0_73849, Y => 
        HIEFFPLA_NET_0_73826);
    
    HIEFFPLA_INST_0_62412 : XA1C
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[1]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73988);
    
    HIEFFPLA_INST_0_65722 : AND3C
      port map(A => HIEFFPLA_NET_0_73298, B => 
        \Science_0/ADC_READ_0/cnt[3]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73299);
    
    HIEFFPLA_INST_0_60075 : MX2
      port map(A => \Science_0_chan5_data[0]\, B => 
        \Science_0_chan5_data[4]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74465);
    
    HIEFFPLA_INST_0_63686 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[1]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_nof_steps[1]_net_1\, S
         => \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73728);
    
    HIEFFPLA_INST_0_64837 : OR3A
      port map(A => HIEFFPLA_NET_0_73528, B => 
        HIEFFPLA_NET_0_73600, C => HIEFFPLA_NET_0_73610, Y => 
        HIEFFPLA_NET_0_73527);
    
    HIEFFPLA_INST_0_66005 : NAND2B
      port map(A => \Science_0/ADC_READ_0/state[0]_net_1\, B => 
        \Science_0/ADC_READ_0/countere\, Y => 
        HIEFFPLA_NET_0_73240);
    
    HIEFFPLA_INST_0_63283 : AND2
      port map(A => \General_Controller_0/uc_rx_state_0[3]_net_1\, 
        B => \General_Controller_0/uc_rx_substate[3]_net_1\, Y
         => HIEFFPLA_NET_0_73789);
    
    HIEFFPLA_INST_0_60464 : MX2
      port map(A => \Science_0_chan4_data[5]\, B => 
        \Science_0_chan4_data[9]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74411);
    
    AFLSDF_INV_32 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_32\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_72697, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\);
    
    \Science_0/ADC_READ_0/cnt2dn[7]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73368, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2dn[7]_net_1\);
    
    \TOP_UART_TX_pad/U0/U0\ : IOPAD_TRI
      port map(D => \TOP_UART_TX_pad/U0/NET1\, E => 
        \TOP_UART_TX_pad/U0/NET2\, PAD => TOP_UART_TX);
    
    HIEFFPLA_INST_0_59131 : NOR3B
      port map(A => HIEFFPLA_NET_0_74719, B => 
        \GS_Readout_0/prevState[3]_net_1\, C => 
        \GS_Readout_0/prevState[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74605);
    
    HIEFFPLA_INST_0_65261 : NOR3A
      port map(A => HIEFFPLA_NET_0_73434, B => 
        \Sensors_0_pressure_raw[11]\, C => 
        \Sensors_0_pressure_raw[18]\, Y => HIEFFPLA_NET_0_73432);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_full\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75367, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/full\);
    
    HIEFFPLA_INST_0_58915 : NOR3B
      port map(A => HIEFFPLA_NET_0_74372, B => 
        HIEFFPLA_NET_0_74371, C => HIEFFPLA_NET_0_74671, Y => 
        HIEFFPLA_NET_0_74660);
    
    \Communications_0/FFU_Command_Checker_0/command_rdy\ : 
        DFN1E0C1
      port map(D => \AFLSDF_INV_27\, CLK => CLKINT_0_Y_0, CLR => 
        CLKINT_1_Y, E => HIEFFPLA_NET_0_75627, Q => 
        Communications_0_ext_rx_rdy);
    
    AFLSDF_INV_2 : INV
      port map(A => \Data_Saving_0/FPGA_Buffer_0/MEMRENEG\, Y => 
        \AFLSDF_INV_2\);
    
    HIEFFPLA_INST_0_66468 : AO1
      port map(A => HIEFFPLA_NET_0_73111, B => 
        HIEFFPLA_NET_0_73132, C => HIEFFPLA_NET_0_73106, Y => 
        HIEFFPLA_NET_0_73112);
    
    HIEFFPLA_INST_0_57261 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[48]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75106);
    
    HIEFFPLA_INST_0_57180 : AO1
      port map(A => \Sensors_0_pressure_time[21]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75082, Y => HIEFFPLA_NET_0_75138);
    
    AFLSDF_INV_8 : INV
      port map(A => Sensors_0_acc_new_data, Y => \AFLSDF_INV_8\);
    
    HIEFFPLA_INST_0_61006 : AOI1B
      port map(A => Eject_Signal_Debounce_0_ffu_ejected_out, B
         => \General_Controller_0/flight_state[2]_net_1\, C => 
        HIEFFPLA_NET_0_74296, Y => HIEFFPLA_NET_0_74298);
    
    HIEFFPLA_INST_0_58517 : NOR3B
      port map(A => HIEFFPLA_NET_0_74738, B => 
        HIEFFPLA_NET_0_74728, C => HIEFFPLA_NET_0_74740, Y => 
        HIEFFPLA_NET_0_74744);
    
    \Communications_0/UART_0/tx_clk_count[2]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75524, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_clk_count_i_0[2]\);
    
    HIEFFPLA_INST_0_63204 : AND3A
      port map(A => HIEFFPLA_NET_0_74118, B => 
        HIEFFPLA_NET_0_74073, C => HIEFFPLA_NET_0_73807, Y => 
        HIEFFPLA_NET_0_73808);
    
    HIEFFPLA_INST_0_58745 : NOR3B
      port map(A => HIEFFPLA_NET_0_74490, B => 
        \GS_Readout_0/state[4]_net_1\, C => HIEFFPLA_NET_0_74725, 
        Y => HIEFFPLA_NET_0_74694);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[7]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[7]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[7]\);
    
    HIEFFPLA_INST_0_57487 : AO1
      port map(A => \Sensors_0_acc_z[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74859, Y => HIEFFPLA_NET_0_75032);
    
    HIEFFPLA_INST_0_59045 : NOR3A
      port map(A => HIEFFPLA_NET_0_74408, B => 
        \GS_Readout_0/state[7]_net_1\, C => HIEFFPLA_NET_0_74643, 
        Y => HIEFFPLA_NET_0_74628);
    
    \Communications_0/UART_0/tx_byte[5]\ : DFN1E1
      port map(D => \GS_Readout_0_send[5]\, CLK => CLKINT_0_Y_0, 
        E => HIEFFPLA_NET_0_75504, Q => 
        \Communications_0/UART_0/tx_byte[5]_net_1\);
    
    HIEFFPLA_INST_0_64616 : NOR3A
      port map(A => HIEFFPLA_NET_0_73619, B => 
        \General_Controller_0/uc_tx_state[1]_net_1\, C => 
        \General_Controller_0/uc_tx_state[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73585);
    
    HIEFFPLA_INST_0_64193 : NOR3A
      port map(A => HIEFFPLA_NET_0_73748, B => 
        \General_Controller_0/uc_tx_state[12]_net_1\, C => 
        \General_Controller_0/uc_tx_state[14]_net_1\, Y => 
        HIEFFPLA_NET_0_73652);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_8\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[1]\\\\\, CLK => 
        CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_8_Q\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[5]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75262, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\);
    
    HIEFFPLA_INST_0_71208 : AOI1A
      port map(A => \Communications_0/UART_1/rx_state[1]_net_1\, 
        B => HIEFFPLA_NET_0_75442, C => HIEFFPLA_NET_0_71973, Y
         => HIEFFPLA_NET_0_75450);
    
    HIEFFPLA_INST_0_70346 : AOI1D
      port map(A => General_Controller_0_st_ren1, B => 
        \SweepTable_0/WEBP\, C => 
        \General_Controller_0_st_raddr_1[5]\, Y => 
        \TableSelect_0_RADDR[5]\);
    
    HIEFFPLA_INST_0_66047 : NOR3B
      port map(A => HIEFFPLA_NET_0_73224, B => 
        \Science_0/DAC_SET_0/state[3]_net_1\, C => 
        HIEFFPLA_NET_0_73223, Y => HIEFFPLA_NET_0_73226);
    
    HIEFFPLA_INST_0_57571 : AO1
      port map(A => \Sensors_0_pressure_raw[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_75004, Y => HIEFFPLA_NET_0_75005);
    
    HIEFFPLA_INST_0_57183 : AO1
      port map(A => \Sensors_0_gyro_time[22]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75136, Y => HIEFFPLA_NET_0_75137);
    
    \Science_0/ADC_READ_0/exp_packet_1[61]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[5]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[61]\);
    
    HIEFFPLA_INST_0_64766 : AND2B
      port map(A => Communications_0_uc_tx_rdy, B => 
        HIEFFPLA_NET_0_73555, Y => HIEFFPLA_NET_0_73546);
    
    \General_Controller_0/sweep_table_samples_per_step[4]\ : 
        DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[4]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[4]_net_1\);
    
    \Communications_0/UART_0/rx_state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75548, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/rx_state[1]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72211, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]_net_1\);
    
    \Science_0/ADC_READ_0/cnt[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73291, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73242, Q => 
        \Science_0/ADC_READ_0/cnt[1]_net_1\);
    
    HIEFFPLA_INST_0_60850 : NAND3C
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, C => 
        \GS_Readout_0/subState[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74343);
    
    \Communications_0/UART_1/rx_clk_count[24]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75464, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75443, Q => 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\);
    
    AFLSDF_INV_0 : INV
      port map(A => \Data_Saving_0/FPGA_Buffer_0/MEMRENEG\, Y => 
        \AFLSDF_INV_0\);
    
    HIEFFPLA_INST_0_70041 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[2]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72237);
    
    HIEFFPLA_INST_0_66012 : AND3
      port map(A => HIEFFPLA_NET_0_73299, B => 
        HIEFFPLA_NET_0_73295, C => 
        \Science_0/ADC_READ_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73238);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[10]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72753, Q => 
        \Sensors_0_acc_z[10]\);
    
    HIEFFPLA_INST_0_68509 : OR3B
      port map(A => GYRO_SCL_c, B => HIEFFPLA_NET_0_72616, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_72633);
    
    \ACCE_SDA_pad/U0/U0\ : IOPAD_BI
      port map(D => \ACCE_SDA_pad/U0/NET1\, E => 
        \ACCE_SDA_pad/U0/NET2\, Y => \ACCE_SDA_pad/U0/NET3\, PAD
         => ACCE_SDA);
    
    \General_Controller_0/gs_id[2]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73922, Q => 
        \General_Controller_0_gs_id[2]\);
    
    \General_Controller_0/uc_rx_state[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73895, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_state[3]_net_1\);
    
    HIEFFPLA_INST_0_66127 : MX2B
      port map(A => \Science_0/DAC_SET_0/vector[11]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73201);
    
    HIEFFPLA_INST_0_61693 : MX2
      port map(A => \SweepTable_0_RD[5]\, B => 
        \SweepTable_1_RD[5]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74159);
    
    HIEFFPLA_INST_0_56374 : AX1D
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, B
         => HIEFFPLA_NET_0_75349, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\, Y
         => HIEFFPLA_NET_0_75297);
    
    \General_Controller_0/sweep_table_step_id[0]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73926, Q => 
        \General_Controller_0/sweep_table_step_id[0]_net_1\);
    
    HIEFFPLA_INST_0_67815 : AO1A
      port map(A => HIEFFPLA_NET_0_72763, B => 
        HIEFFPLA_NET_0_72771, C => HIEFFPLA_NET_0_72794, Y => 
        HIEFFPLA_NET_0_72795);
    
    \Science_0/ADC_READ_0/cnt3up[4]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73332, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3up[4]_net_1\);
    
    \Science_0/SET_LP_GAIN_0/state[6]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73153, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/state[6]_net_1\);
    
    HIEFFPLA_INST_0_69336 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72415);
    
    \General_Controller_0/status_new_data\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74267, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        General_Controller_0_status_new_data);
    
    \Science_0/ADC_READ_0/chan3_data[11]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[17]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[11]\);
    
    HIEFFPLA_INST_0_67739 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, B
         => HIEFFPLA_NET_0_72935, Y => HIEFFPLA_NET_0_72812);
    
    HIEFFPLA_INST_0_65783 : AND3
      port map(A => HIEFFPLA_NET_0_73238, B => 
        \Science_0/ADC_READ_0/cnt_chan[0]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt_chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73280);
    
    HIEFFPLA_INST_0_57483 : AO1
      port map(A => \Sensors_0_acc_z[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74861, Y => HIEFFPLA_NET_0_75033);
    
    \Science_0/ADC_READ_0/exp_packet_1[29]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[13]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[29]\);
    
    \Communications_0/UART_1/tx_rdy\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75386, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => Communications_0_uc_tx_rdy);
    
    HIEFFPLA_INST_0_59330 : MX2
      port map(A => \Science_0_chan4_data[7]\, B => 
        \Science_0_chan4_data[11]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74567);
    
    \General_Controller_0/state_seconds[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74240, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[0]_net_1\);
    
    HIEFFPLA_INST_0_54959 : AO1A
      port map(A => General_Controller_0_ext_oen, B => 
        \Communications_0/FFU_Command_Checker_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_75626, Y => HIEFFPLA_NET_0_75627);
    
    \Data_Saving_0/Packet_Saver_0/old_mag_new_data\ : DFN0P1
      port map(D => \AFLSDF_INV_28\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => 
        \Data_Saving_0/Packet_Saver_0/old_mag_new_data_i_0\);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72340, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[0]_net_1\);
    
    HIEFFPLA_INST_0_66828 : AO1
      port map(A => HIEFFPLA_NET_0_73019, B => 
        HIEFFPLA_NET_0_73055, C => HIEFFPLA_NET_0_73016, Y => 
        HIEFFPLA_NET_0_73026);
    
    HIEFFPLA_INST_0_66528 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[3]_net_1\, 
        B => ACCE_SCL_c, C => HIEFFPLA_NET_0_73143, Y => 
        HIEFFPLA_NET_0_73101);
    
    \Communications_0/UART_1/rx_byte[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75378, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75494, Q => 
        \Communications_0/UART_1/rx_byte[2]_net_1\);
    
    HIEFFPLA_INST_0_56758 : AOI1B
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[1]_net_1\, B => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_75179, Y => HIEFFPLA_NET_0_75214);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_5\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[2]\\\\\, CLK => 
        CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_5_Q\);
    
    \AB_pad/U0/U1\ : IOIN_IB
      port map(YIN => \AB_pad/U0/NET1\, Y => AB_c);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRY[2]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75303, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[2]\\\\\);
    
    \Science_0/ADC_READ_0/cnt2dn[2]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73374, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2dn[2]_net_1\);
    
    HIEFFPLA_INST_0_60741 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[40]\, B => 
        \Data_Hub_Packets_0_status_packet[44]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74365);
    
    HIEFFPLA_INST_0_56652 : MX2
      port map(A => HIEFFPLA_NET_0_75195, B => 
        HIEFFPLA_NET_0_75061, S => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75228);
    
    HIEFFPLA_INST_0_67172 : AND3
      port map(A => HIEFFPLA_NET_0_72959, B => 
        HIEFFPLA_NET_0_72956, C => HIEFFPLA_NET_0_72950, Y => 
        HIEFFPLA_NET_0_72946);
    
    HIEFFPLA_INST_0_57012 : MX2
      port map(A => HIEFFPLA_NET_0_75042, B => 
        HIEFFPLA_NET_0_74958, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75182);
    
    \General_Controller_0/sweep_table_nof_steps[2]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73980, Q => 
        \General_Controller_0/sweep_table_nof_steps[2]_net_1\);
    
    \ACST_pad/U0/U0\ : IOPAD_TRI
      port map(D => \ACST_pad/U0/NET1\, E => \ACST_pad/U0/NET2\, 
        PAD => ACST);
    
    HIEFFPLA_INST_0_67130 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[7]_net_1\, 
        B => HIEFFPLA_NET_0_72879, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72958);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72356, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_net_1\);
    
    HIEFFPLA_INST_0_61765 : XOR2
      port map(A => HIEFFPLA_NET_0_74149, B => 
        \General_Controller_0/sweep_table_sweep_cnt[11]_net_1\, Y
         => HIEFFPLA_NET_0_74142);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/data_out[0]\ : 
        DFN0E1C1
      port map(D => ACCE_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73125, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\);
    
    HIEFFPLA_INST_0_55883 : AO1D
      port map(A => HIEFFPLA_NET_0_75420, B => 
        HIEFFPLA_NET_0_75386, C => HIEFFPLA_NET_0_75404, Y => 
        HIEFFPLA_NET_0_75405);
    
    \Timekeeper_0/milliseconds[22]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72102, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[22]\);
    
    HIEFFPLA_INST_0_65273 : NOR2A
      port map(A => HIEFFPLA_NET_0_73468, B => 
        \Sensors_0_pressure_raw[14]\, Y => HIEFFPLA_NET_0_73428);
    
    HIEFFPLA_INST_0_64277 : MX2
      port map(A => HIEFFPLA_NET_0_73738, B => 
        HIEFFPLA_NET_0_73730, S => HIEFFPLA_NET_0_73588, Y => 
        HIEFFPLA_NET_0_73642);
    
    HIEFFPLA_INST_0_59246 : NOR3B
      port map(A => \GS_Readout_0/subState[1]_net_1\, B => 
        HIEFFPLA_NET_0_74634, C => \GS_Readout_0/state[6]_net_1\, 
        Y => HIEFFPLA_NET_0_74580);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72868, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_68342 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, B => 
        HIEFFPLA_NET_0_72676, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_72677);
    
    HIEFFPLA_INST_0_61813 : AND2
      port map(A => 
        \General_Controller_0/sweep_table_write_wait[0]_net_1\, B
         => 
        \General_Controller_0/sweep_table_write_wait[1]_net_1\, Y
         => HIEFFPLA_NET_0_74124);
    
    HIEFFPLA_INST_0_61248 : XA1C
      port map(A => HIEFFPLA_NET_0_74251, B => 
        \General_Controller_0/state_seconds[12]_net_1\, C => 
        HIEFFPLA_NET_0_74217, Y => HIEFFPLA_NET_0_74237);
    
    HIEFFPLA_INST_0_70727 : AND3
      port map(A => \Timing_0/m_count[3]_net_1\, B => 
        \Timing_0/m_count[4]_net_1\, C => 
        \Timing_0/m_count[5]_net_1\, Y => HIEFFPLA_NET_0_72030);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[8]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[8]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[8]\);
    
    HIEFFPLA_INST_0_55235 : MX2A
      port map(A => HIEFFPLA_NET_0_75594, B => 
        HIEFFPLA_NET_0_75545, S => 
        \Communications_0/UART_0/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75555);
    
    HIEFFPLA_INST_0_57396 : AO1
      port map(A => \Science_0_exp_packet_0[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74851, Y => HIEFFPLA_NET_0_75057);
    
    HIEFFPLA_INST_0_68552 : AO1
      port map(A => HIEFFPLA_NET_0_72620, B => GYRO_SCL_c, C => 
        HIEFFPLA_NET_0_72621, Y => HIEFFPLA_NET_0_72619);
    
    HIEFFPLA_INST_0_67887 : AOI1
      port map(A => HIEFFPLA_NET_0_72940, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        C => HIEFFPLA_NET_0_72779, Y => HIEFFPLA_NET_0_72780);
    
    HIEFFPLA_INST_0_61136 : AO1
      port map(A => \s_clks_net_0[24]\, B => 
        \General_Controller_0/old_1Hz_i_0\, C => 
        HIEFFPLA_NET_0_74217, Y => HIEFFPLA_NET_0_74268);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[8]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_75245, CLK => CLKINT_0_Y_0, E
         => CLKINT_1_Y, Q => 
        \Data_Saving_0/Interrupt_Generator_0/counter[8]_net_1\);
    
    \Science_0/SET_LP_GAIN_0/L1WR\ : DFN0C1
      port map(D => \Science_0/SET_LP_GAIN_0/state_i_0[3]\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => L1WR_c);
    
    \PRESSURE_SDA_pad/U0/U1\ : IOBI_IB_OB_EB
      port map(D => 
        \Sensors_0.Pressure_Sensor_0.I2C_Master_0.sda_1\, E => 
        sda_cl_1_RNIGPAD, YIN => \PRESSURE_SDA_pad/U0/NET3\, DOUT
         => \PRESSURE_SDA_pad/U0/NET1\, EOUT => 
        \PRESSURE_SDA_pad/U0/NET2\, Y => PRESSURE_SDA_in);
    
    HIEFFPLA_INST_0_70944 : NAND3C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72003);
    
    \FMC_NOE_pad/U0/U0\ : IOPAD_IN
      port map(PAD => FMC_NOE, Y => \FMC_NOE_pad/U0/NET1\);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_18\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[5]\\\\\, CLK => 
        CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_18_Q\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/data_out_rdy\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72699, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72672, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\);
    
    HIEFFPLA_INST_0_62918 : NOR3B
      port map(A => HIEFFPLA_NET_0_73908, B => 
        Communications_0_uc_rx_rdy, C => HIEFFPLA_NET_0_73889, Y
         => HIEFFPLA_NET_0_73866);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[1]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72276, Q => \Sensors_0_pressure_raw[1]\);
    
    HIEFFPLA_INST_0_67256 : AO1
      port map(A => HIEFFPLA_NET_0_72784, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_72925, Y => HIEFFPLA_NET_0_72926);
    
    HIEFFPLA_INST_0_56712 : MX2
      port map(A => HIEFFPLA_NET_0_75189, B => 
        HIEFFPLA_NET_0_75049, S => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75222);
    
    \General_Controller_0/uc_oen\ : DFN1E0C1
      port map(D => Communications_0_uc_rx_rdy, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74121, Q => General_Controller_0_uc_oen);
    
    HIEFFPLA_INST_0_69465 : OR2A
      port map(A => HIEFFPLA_NET_0_72381, B => 
        HIEFFPLA_NET_0_72392, Y => HIEFFPLA_NET_0_72382);
    
    HIEFFPLA_INST_0_58736 : NOR3B
      port map(A => HIEFFPLA_NET_0_74627, B => 
        HIEFFPLA_NET_0_74386, C => HIEFFPLA_NET_0_74510, Y => 
        HIEFFPLA_NET_0_74695);
    
    \Communications_0/UART_1/tx_count[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75392, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75388, Q => 
        \Communications_0/UART_1/tx_count[1]_net_1\);
    
    \General_Controller_0/st_wdata[2]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[2]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[2]\);
    
    HIEFFPLA_INST_0_69267 : OR3A
      port map(A => HIEFFPLA_NET_0_72491, B => 
        HIEFFPLA_NET_0_72431, C => HIEFFPLA_NET_0_72499, Y => 
        HIEFFPLA_NET_0_72433);
    
    HIEFFPLA_INST_0_67695 : AO1
      port map(A => HIEFFPLA_NET_0_72812, B => 
        HIEFFPLA_NET_0_72811, C => HIEFFPLA_NET_0_72847, Y => 
        HIEFFPLA_NET_0_72822);
    
    HIEFFPLA_INST_0_57502 : AOI1
      port map(A => \Science_0_exp_packet_0[20]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_75026, Y => HIEFFPLA_NET_0_75027);
    
    \General_Controller_0/st_wdata[3]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[3]\);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_0[8]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74766, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[1]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[1]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[1]\);
    
    HIEFFPLA_INST_0_66255 : XOR2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G4[0]_net_1\, B
         => \Science_0/ADC_READ_0_G4[0]\, Y => 
        HIEFFPLA_NET_0_73165);
    
    HIEFFPLA_INST_0_70956 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[0]\, 
        C => HIEFFPLA_NET_0_72978, Y => HIEFFPLA_NET_0_72001);
    
    HIEFFPLA_INST_0_57108 : MX2
      port map(A => HIEFFPLA_NET_0_74935, B => 
        HIEFFPLA_NET_0_74878, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75166);
    
    \Science_0/ADC_READ_0/chan5_data[11]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[17]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[11]\);
    
    HIEFFPLA_INST_0_67230 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_72761, Y => HIEFFPLA_NET_0_72933);
    
    HIEFFPLA_INST_0_59088 : AND2
      port map(A => General_Controller_0_readout_en, B => 
        \GS_Readout_0/state[7]_net_1\, Y => HIEFFPLA_NET_0_74616);
    
    HIEFFPLA_INST_0_69308 : NOR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\, 
        B => HIEFFPLA_NET_0_72350, C => HIEFFPLA_NET_0_72427, Y
         => HIEFFPLA_NET_0_72422);
    
    HIEFFPLA_INST_0_66199 : AO1
      port map(A => \Science_0/SET_LP_GAIN_0/state[4]_net_1\, B
         => \Science_0/ADC_READ_0_G4[1]\, C => 
        HIEFFPLA_NET_0_73167, Y => HIEFFPLA_NET_0_73180);
    
    HIEFFPLA_INST_0_64775 : AOI1C
      port map(A => HIEFFPLA_NET_0_73605, B => 
        HIEFFPLA_NET_0_73541, C => 
        \General_Controller_0/uc_tx_state[14]_net_1\, Y => 
        HIEFFPLA_NET_0_73543);
    
    HIEFFPLA_INST_0_62638 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[3]_net_1\, 
        B => \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        HIEFFPLA_NET_0_73909, Y => HIEFFPLA_NET_0_73940);
    
    HIEFFPLA_INST_0_61657 : MX2
      port map(A => \SweepTable_0_RD[14]\, B => 
        \SweepTable_1_RD[14]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74165);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[0]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72503, Q => 
        \Sensors_0_gyro_x[0]\);
    
    HIEFFPLA_INST_0_66768 : AO1
      port map(A => HIEFFPLA_NET_0_73052, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        C => HIEFFPLA_NET_0_73099, Y => HIEFFPLA_NET_0_73039);
    
    \General_Controller_0/sweep_table_probe_id[6]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73924, Q => 
        \General_Controller_0/sweep_table_probe_id[6]_net_1\);
    
    HIEFFPLA_INST_0_58242 : AO1
      port map(A => \Sensors_0_gyro_time[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75114, Y => HIEFFPLA_NET_0_74822);
    
    \Science_0/ADC_READ_0/chan2_data[4]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[4]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[2]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72503, Q => 
        \Sensors_0_gyro_x[2]\);
    
    \General_Controller_0/sweep_table_write_wait[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74122, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/sweep_table_write_wait[1]_net_1\);
    
    HIEFFPLA_INST_0_68471 : OR3B
      port map(A => HIEFFPLA_NET_0_72640, B => 
        HIEFFPLA_NET_0_72642, C => \Sensors_0/Gyro_0/state[8]\, Y
         => HIEFFPLA_NET_0_72643);
    
    HIEFFPLA_INST_0_67460 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        B => HIEFFPLA_NET_0_72717, C => HIEFFPLA_NET_0_72744, Y
         => HIEFFPLA_NET_0_72873);
    
    HIEFFPLA_INST_0_67721 : NOR2A
      port map(A => HIEFFPLA_NET_0_72844, B => 
        HIEFFPLA_NET_0_72798, Y => HIEFFPLA_NET_0_72816);
    
    HIEFFPLA_INST_0_57441 : AO1B
      port map(A => \Sensors_0_mag_z[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75044, Y => HIEFFPLA_NET_0_75045);
    
    \Timekeeper_0/milliseconds[11]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72114, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[11]\);
    
    HIEFFPLA_INST_0_58798 : NOR3A
      port map(A => HIEFFPLA_NET_0_74667, B => 
        HIEFFPLA_NET_0_74670, C => HIEFFPLA_NET_0_74699, Y => 
        HIEFFPLA_NET_0_74682);
    
    \Communications_0/UART_1/rx_clk_count[26]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75461, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75443, Q => 
        \Communications_0/UART_1/rx_clk_count[26]_net_1\);
    
    HIEFFPLA_INST_0_64986 : AO1B
      port map(A => HIEFFPLA_NET_0_73483, B => 
        HIEFFPLA_NET_0_73482, C => HIEFFPLA_NET_0_73477, Y => 
        HIEFFPLA_NET_0_73495);
    
    HIEFFPLA_INST_0_60797 : MX2
      port map(A => HIEFFPLA_NET_0_74444, B => 
        HIEFFPLA_NET_0_74440, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74357);
    
    HIEFFPLA_INST_0_67994 : AND3C
      port map(A => HIEFFPLA_NET_0_72739, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72759);
    
    HIEFFPLA_INST_0_61222 : NAND2
      port map(A => \General_Controller_0/state_seconds[6]_net_1\, 
        B => \General_Controller_0/state_seconds[5]_net_1\, Y => 
        HIEFFPLA_NET_0_74245);
    
    HIEFFPLA_INST_0_59166 : NAND3A
      port map(A => \GS_Readout_0/prevState[7]_net_1\, B => 
        HIEFFPLA_NET_0_74724, C => HIEFFPLA_NET_0_74720, Y => 
        HIEFFPLA_NET_0_74597);
    
    HIEFFPLA_INST_0_55783 : MX2
      port map(A => HIEFFPLA_NET_0_75424, B => 
        HIEFFPLA_NET_0_75423, S => 
        \Communications_0/UART_1/tx_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75426);
    
    HIEFFPLA_INST_0_67562 : AO1
      port map(A => HIEFFPLA_NET_0_72947, B => 
        HIEFFPLA_NET_0_72957, C => HIEFFPLA_NET_0_72825, Y => 
        HIEFFPLA_NET_0_72851);
    
    HIEFFPLA_INST_0_65443 : XA1C
      port map(A => \Science_0/ADC_READ_0/cnt2dn[2]_net_1\, B => 
        HIEFFPLA_NET_0_73380, C => HIEFFPLA_NET_0_73381, Y => 
        HIEFFPLA_NET_0_73374);
    
    HIEFFPLA_INST_0_70517 : AX1C
      port map(A => \Timekeeper_0_milliseconds[1]\, B => 
        \Timekeeper_0_milliseconds[0]\, C => 
        \Timekeeper_0_milliseconds[2]\, Y => HIEFFPLA_NET_0_72100);
    
    HIEFFPLA_INST_0_68181 : AX1
      port map(A => HIEFFPLA_NET_0_72764, B => 
        HIEFFPLA_NET_0_72716, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72713);
    
    HIEFFPLA_INST_0_66166 : MX2B
      port map(A => \Science_0/DAC_SET_0/vector[3]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73192);
    
    HIEFFPLA_INST_0_59261 : XA1
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, C => 
        HIEFFPLA_NET_0_74544, Y => HIEFFPLA_NET_0_74578);
    
    \General_Controller_0/sweep_table_points[13]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[13]_net_1\);
    
    HIEFFPLA_INST_0_58141 : AO1
      port map(A => \Sensors_0_mag_time[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75148, Y => HIEFFPLA_NET_0_74841);
    
    \Science_0/ADC_READ_0/exp_packet_1[0]\ : DFN1E0
      port map(D => \AFLSDF_INV_29\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[0]\);
    
    HIEFFPLA_INST_0_59848 : MX2
      port map(A => \Sensors_0_pressure_temp_raw[14]\, B => 
        \Sensors_0_pressure_temp_raw[18]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74498);
    
    \Science_0/ADC_READ_0/g3i[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73254, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73419, Q => 
        \Science_0/ADC_READ_0_G3[1]\);
    
    HIEFFPLA_INST_0_61798 : NOR2A
      port map(A => HIEFFPLA_NET_0_73918, B => 
        HIEFFPLA_NET_0_74126, Y => HIEFFPLA_NET_0_74127);
    
    HIEFFPLA_INST_0_54967 : NOR2A
      port map(A => \Communications_0/UART_0_rx_rdy\, B => 
        \Communications_0/FFU_Command_Checker_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_75624);
    
    HIEFFPLA_INST_0_70671 : XOR2
      port map(A => \s_time[5]\, B => HIEFFPLA_NET_0_72038, Y => 
        HIEFFPLA_NET_0_72049);
    
    HIEFFPLA_INST_0_62436 : AOI1
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state[3]_net_1\, C => 
        HIEFFPLA_NET_0_73982, Y => HIEFFPLA_NET_0_73983);
    
    \Science_0/ADC_READ_0/data_b[15]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[15]_net_1\);
    
    HIEFFPLA_INST_0_70533 : NOR2A
      port map(A => \m_time[7]\, B => 
        \Timekeeper_0/old_1kHz_net_1\, Y => HIEFFPLA_NET_0_72091);
    
    HIEFFPLA_INST_0_66139 : MX2
      port map(A => \Science_0/DAC_SET_0/vector[15]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[0]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73197);
    
    \Data_Saving_0/Packet_Saver_0/old_status_new_data\ : DFN0P1
      port map(D => \AFLSDF_INV_30\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => 
        \Data_Saving_0/Packet_Saver_0/old_status_new_data_i_0\);
    
    HIEFFPLA_INST_0_58469 : NOR2A
      port map(A => HIEFFPLA_NET_0_74766, B => 
        \Data_Saving_0/Packet_Saver_0/status_flag_net_1\, Y => 
        HIEFFPLA_NET_0_74759);
    
    \Sensors_0/Gyro_0/I2C_Master_0/state[8]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_72604, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/state[8]\);
    
    HIEFFPLA_INST_0_63866 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[7]_net_1\, B
         => 
        \General_Controller_0/sweep_table_sample_skip[7]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73698);
    
    HIEFFPLA_INST_0_61986 : AND2B
      port map(A => \General_Controller_0/uc_rx_byte[3]_net_1\, B
         => \General_Controller_0/uc_rx_byte[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74081);
    
    HIEFFPLA_INST_0_58375 : AND2
      port map(A => \Sensors_0_mag_z[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        Y => HIEFFPLA_NET_0_74787);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_9\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[2]\\\\\, CLK => 
        CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_9_Q\);
    
    \Science_0/DAC_SET_0/vector[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73195, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[1]_net_1\);
    
    HIEFFPLA_INST_0_62143 : NAND3C
      port map(A => HIEFFPLA_NET_0_74032, B => 
        HIEFFPLA_NET_0_73945, C => HIEFFPLA_NET_0_73996, Y => 
        HIEFFPLA_NET_0_74043);
    
    HIEFFPLA_INST_0_70765 : XA1C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[0]_net_1\, 
        B => \Sensors_0/Pressure_Sensor_0/state[8]\, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72018);
    
    HIEFFPLA_INST_0_65693 : NAND2B
      port map(A => CLKINT_1_Y, B => 
        \Science_0/ADC_READ_0/cnt4up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73308);
    
    HIEFFPLA_INST_0_62904 : NAND2A
      port map(A => \General_Controller_0/uc_rx_state[4]_net_1\, 
        B => \General_Controller_0/uc_rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73869);
    
    HIEFFPLA_INST_0_57188 : AO1
      port map(A => \Sensors_0_pressure_time[23]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75081, Y => HIEFFPLA_NET_0_75135);
    
    HIEFFPLA_INST_0_55518 : NOR3B
      port map(A => HIEFFPLA_NET_0_75452, B => 
        HIEFFPLA_NET_0_75488, C => 
        \Communications_0/UART_1/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75490);
    
    HIEFFPLA_INST_0_62559 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state[3]_net_1\, 
        B => \General_Controller_0/uc_rx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_73909, Y => HIEFFPLA_NET_0_73957);
    
    \General_Controller_0/sweep_table_sweep_cnt[11]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74142, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[11]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[15]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72283, Q => 
        \Sensors_0_pressure_temp_raw[15]\);
    
    \PRESSURE_SDA_pad/U0/U0\ : IOPAD_BI
      port map(D => \PRESSURE_SDA_pad/U0/NET1\, E => 
        \PRESSURE_SDA_pad/U0/NET2\, Y => 
        \PRESSURE_SDA_pad/U0/NET3\, PAD => PRESSURE_SDA);
    
    HIEFFPLA_INST_0_56389 : AND3A
      port map(A => \Data_Saving_0/FPGA_Buffer_0/full\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[0]\\\\\, C
         => \Data_Saving_0/Packet_Saver_0_we\, Y => 
        HIEFFPLA_NET_0_75293);
    
    \Science_0/ADC_READ_0/data_b[6]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[5]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[6]_net_1\);
    
    HIEFFPLA_INST_0_66553 : AO1
      port map(A => HIEFFPLA_NET_0_73091, B => 
        \Sensors_0.Accelerometer_0.I2C_Master_0.sda_1\, C => 
        HIEFFPLA_NET_0_73083, Y => HIEFFPLA_NET_0_73093);
    
    HIEFFPLA_INST_0_65546 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt3dn[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt3dn[0]_net_1\, C => 
        HIEFFPLA_NET_0_73349, Y => HIEFFPLA_NET_0_73346);
    
    HIEFFPLA_INST_0_63218 : NAND2B
      port map(A => 
        \General_Controller_0/uc_rx_substate[4]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73804);
    
    HIEFFPLA_INST_0_55821 : AO1
      port map(A => HIEFFPLA_NET_0_75415, B => 
        HIEFFPLA_NET_0_75413, C => 
        \Communications_0/UART_1/tx_clk_count_i_0[8]\, Y => 
        HIEFFPLA_NET_0_75420);
    
    HIEFFPLA_INST_0_68295 : AX1B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_72684, Y => HIEFFPLA_NET_0_72687);
    
    HIEFFPLA_INST_0_56987 : AOI1C
      port map(A => HIEFFPLA_NET_0_74891, B => 
        HIEFFPLA_NET_0_75047, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75186);
    
    HIEFFPLA_INST_0_56232 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, B
         => HIEFFPLA_NET_0_75370, C => HIEFFPLA_NET_0_75273, Y
         => HIEFFPLA_NET_0_75329);
    
    HIEFFPLA_INST_0_71004 : AOI1
      port map(A => HIEFFPLA_NET_0_71993, B => 
        HIEFFPLA_NET_0_73473, C => HIEFFPLA_NET_0_73497, Y => 
        HIEFFPLA_NET_0_73475);
    
    HIEFFPLA_INST_0_58402 : AO1
      port map(A => \Sensors_0_pressure_raw[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74777, Y => HIEFFPLA_NET_0_74778);
    
    HIEFFPLA_INST_0_63416 : MX2
      port map(A => HIEFFPLA_NET_0_73757, B => 
        HIEFFPLA_NET_0_73691, S => HIEFFPLA_NET_0_73608, Y => 
        HIEFFPLA_NET_0_73765);
    
    \Communications_0/UART_1/rx_byte[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75378, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75490, Q => 
        \Communications_0/UART_1/rx_byte[6]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72535, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\);
    
    \Science_0/ADC_READ_0/cnt1dn[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73401, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1dn[7]_net_1\);
    
    HIEFFPLA_INST_0_69224 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, B
         => HIEFFPLA_NET_0_72491, C => HIEFFPLA_NET_0_72540, Y
         => HIEFFPLA_NET_0_72444);
    
    HIEFFPLA_INST_0_60107 : MX2
      port map(A => \Science_0_chan3_data[9]\, B => 
        \Science_0_chan2_data[1]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74461);
    
    HIEFFPLA_INST_0_66618 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]_net_1\, 
        B => ACCE_SCL_c, C => HIEFFPLA_NET_0_73080, Y => 
        HIEFFPLA_NET_0_73081);
    
    HIEFFPLA_INST_0_61217 : OA1C
      port map(A => \General_Controller_0/state_seconds[3]_net_1\, 
        B => HIEFFPLA_NET_0_74263, C => 
        \General_Controller_0/state_seconds[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74247);
    
    HIEFFPLA_INST_0_64501 : AOI1C
      port map(A => HIEFFPLA_NET_0_73586, B => 
        \General_Controller_0/uc_tx_state[3]_net_1\, C => 
        HIEFFPLA_NET_0_73559, Y => HIEFFPLA_NET_0_73613);
    
    HIEFFPLA_INST_0_62350 : NAND3B
      port map(A => HIEFFPLA_NET_0_73977, B => 
        HIEFFPLA_NET_0_74044, C => HIEFFPLA_NET_0_73999, Y => 
        HIEFFPLA_NET_0_74000);
    
    HIEFFPLA_INST_0_55753 : AO1
      port map(A => HIEFFPLA_NET_0_75453, B => 
        HIEFFPLA_NET_0_75430, C => HIEFFPLA_NET_0_75439, Y => 
        HIEFFPLA_NET_0_75432);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/data_out_1[1]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_72569, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72547, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[1]\);
    
    \Science_0/ADC_READ_0/chan6_data[2]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[2]\);
    
    \Science_0/ADC_READ_0/chan0_data[2]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[2]\);
    
    HIEFFPLA_INST_0_58212 : AO1
      port map(A => \Sensors_0_gyro_x[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74826, Y => HIEFFPLA_NET_0_74827);
    
    HIEFFPLA_INST_0_70423 : AX1C
      port map(A => \Timekeeper_0_microseconds[22]\, B => 
        HIEFFPLA_NET_0_72153, C => 
        \Timekeeper_0_microseconds[23]\, Y => 
        HIEFFPLA_NET_0_72136);
    
    HIEFFPLA_INST_0_68346 : NAND3
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, C => 
        GYRO_SCL_c, Y => HIEFFPLA_NET_0_72676);
    
    AFLSDF_INV_6 : INV
      port map(A => CLKINT_1_Y, Y => \AFLSDF_INV_6\);
    
    HIEFFPLA_INST_0_58609 : NOR3A
      port map(A => HIEFFPLA_NET_0_74721, B => 
        \GS_Readout_0/prevState[5]_net_1\, C => 
        \GS_Readout_0/prevState[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74720);
    
    HIEFFPLA_INST_0_56131 : AO13
      port map(A => HIEFFPLA_NET_0_75338, B => 
        HIEFFPLA_NET_0_75315, C => HIEFFPLA_NET_0_75272, Y => 
        HIEFFPLA_NET_0_75340);
    
    HIEFFPLA_INST_0_61460 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[50]\, B => 
        \Timekeeper_0_milliseconds[10]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74196);
    
    \General_Controller_0/unit_id[4]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73990, Q => 
        \General_Controller_0_unit_id[4]\);
    
    HIEFFPLA_INST_0_70461 : AND2
      port map(A => HIEFFPLA_NET_0_72126, B => 
        \Timekeeper_0_milliseconds[21]\, Y => 
        HIEFFPLA_NET_0_72122);
    
    HIEFFPLA_INST_0_65401 : OR2A
      port map(A => \Science_0/ADC_READ_0/cnt2dn[3]_net_1\, B => 
        HIEFFPLA_NET_0_73377, Y => HIEFFPLA_NET_0_73387);
    
    HIEFFPLA_INST_0_68921 : NOR3B
      port map(A => HIEFFPLA_NET_0_72501, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, C
         => \Sensors_0/Gyro_0/I2C_Master_0_s_ack_error\, Y => 
        HIEFFPLA_NET_0_72521);
    
    \General_Controller_0/st_wdata[7]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[7]\);
    
    HIEFFPLA_INST_0_56771 : AOI1C
      port map(A => HIEFFPLA_NET_0_75176, B => 
        HIEFFPLA_NET_0_75177, C => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75212);
    
    HIEFFPLA_INST_0_65967 : AO1A
      port map(A => HIEFFPLA_NET_0_73247, B => 
        HIEFFPLA_NET_0_73245, C => HIEFFPLA_NET_0_73249, Y => 
        HIEFFPLA_NET_0_73250);
    
    \RESET_pad/U0/U0\ : IOPAD_IN
      port map(PAD => RESET, Y => \RESET_pad/U0/NET1\);
    
    HIEFFPLA_INST_0_62649 : AND2
      port map(A => HIEFFPLA_NET_0_73775, B => 
        \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73937);
    
    HIEFFPLA_INST_0_69201 : AO1A
      port map(A => HIEFFPLA_NET_0_72557, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        C => HIEFFPLA_NET_0_72441, Y => HIEFFPLA_NET_0_72448);
    
    HIEFFPLA_INST_0_63716 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[6]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_nof_steps[6]_net_1\, S
         => \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73723);
    
    HIEFFPLA_INST_0_88367 : AO18
      port map(A => HIEFFPLA_NET_0_88384, B => 
        HIEFFPLA_NET_0_89694, C => HIEFFPLA_NET_0_88385, Y => 
        HIEFFPLA_NET_0_88387);
    
    \Communications_0/UART_1/recv[5]\ : DFN1E1C1
      port map(D => \Communications_0/UART_1/rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75441, Q => \Communications_0_uc_recv[5]\);
    
    HIEFFPLA_INST_0_66544 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        B => \Sensors_0/Accelerometer_0/state_0[8]\, Y => 
        HIEFFPLA_NET_0_73095);
    
    \L1WR_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => L1WR_c, E => \VCC\, DOUT => 
        \L1WR_pad/U0/NET1\, EOUT => \L1WR_pad/U0/NET2\);
    
    \General_Controller_0/status_bits_1[37]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74207, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[4]\);
    
    HIEFFPLA_INST_0_65531 : AND3
      port map(A => HIEFFPLA_NET_0_73356, B => 
        HIEFFPLA_NET_0_73353, C => HIEFFPLA_NET_0_73277, Y => 
        HIEFFPLA_NET_0_73350);
    
    HIEFFPLA_INST_0_58111 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_74850);
    
    \General_Controller_0/flight_state[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74289, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/flight_state[3]_net_1\);
    
    HIEFFPLA_INST_0_55926 : AO1D
      port map(A => HIEFFPLA_NET_0_75387, B => 
        \Communications_0/UART_1/tx_count[0]_net_1\, C => 
        HIEFFPLA_NET_0_75396, Y => HIEFFPLA_NET_0_75393);
    
    \Timing_0/s_count[5]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72052, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_count[5]_net_1\);
    
    \UC_I2C4_SCL_pad/U0/U1\ : IOIN_IB
      port map(YIN => \UC_I2C4_SCL_pad/U0/NET1\, Y => 
        FRAM_SCL_c_c);
    
    HIEFFPLA_INST_0_57601 : AO1
      port map(A => \Sensors_0_pressure_raw[13]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74995, Y => HIEFFPLA_NET_0_74996);
    
    \Communications_0/UART_1/tx_byte[5]\ : DFN1E1
      port map(D => \General_Controller_0_uc_send[5]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_75385, Q => 
        \Communications_0/UART_1/tx_byte[5]_net_1\);
    
    \Science_0/ADC_READ_0/chan4_data[1]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[1]\);
    
    HIEFFPLA_INST_0_62523 : OR2A
      port map(A => HIEFFPLA_NET_0_74013, B => 
        HIEFFPLA_NET_0_74015, Y => HIEFFPLA_NET_0_73965);
    
    HIEFFPLA_INST_0_57771 : AO1
      port map(A => \Sensors_0_pressure_raw[19]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, C
         => HIEFFPLA_NET_0_74946, Y => HIEFFPLA_NET_0_74947);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[6]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[6]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[6]\);
    
    \Science_0/ADC_READ_0/chan5_data[3]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[3]\);
    
    \Timekeeper_0/milliseconds[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72096, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[6]\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/scl\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_72633, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        GYRO_SCL_c);
    
    \Timing_0/s_time[8]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72041, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_time[8]_net_1\);
    
    HIEFFPLA_INST_0_55363 : NAND3C
      port map(A => HIEFFPLA_NET_0_75536, B => 
        \Communications_0/UART_0/tx_clk_count_i_0[3]\, C => 
        \Communications_0/UART_0/tx_clk_count_i_0[4]\, Y => 
        HIEFFPLA_NET_0_75529);
    
    HIEFFPLA_INST_0_68467 : AND3
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_net_1\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_1_net_1\, C
         => \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_2_net_1\, Y => 
        sda_cl_1_RNITJT01);
    
    \Science_0/ADC_READ_0/g1i[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73264, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0_G1[1]\);
    
    HIEFFPLA_INST_0_63061 : NOR2A
      port map(A => HIEFFPLA_NET_0_73837, B => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73838);
    
    HIEFFPLA_INST_0_57768 : AOI1
      port map(A => \Sensors_0_gyro_time[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74831, Y => HIEFFPLA_NET_0_74948);
    
    HIEFFPLA_INST_0_55811 : MX2C
      port map(A => \Communications_0/UART_1/tx_byte[1]_net_1\, B
         => \Communications_0/UART_1/tx_byte[5]_net_1\, S => 
        \Communications_0/UART_1/tx_count[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75422);
    
    HIEFFPLA_INST_0_70630 : AND2
      port map(A => \Timing_0/s_count[7]_net_1\, B => 
        \Timing_0/s_count[3]_net_1\, Y => HIEFFPLA_NET_0_72059);
    
    \Communications_0/FFU_Command_Checker_0/command_out[7]\ : 
        DFN1E1C1
      port map(D => \Communications_0/UART_0_recv[7]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75625, Q => \Communications_0_ext_recv[7]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[21]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72280, Q => \Sensors_0_pressure_raw[21]\);
    
    HIEFFPLA_INST_0_64634 : NOR3B
      port map(A => HIEFFPLA_NET_0_73592, B => 
        HIEFFPLA_NET_0_73580, C => 
        \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73581);
    
    HIEFFPLA_INST_0_56418 : MX2
      port map(A => \FMC_DA_c[2]\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[2]\\\\\, S => 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\, Y => 
        HIEFFPLA_NET_0_75285);
    
    HIEFFPLA_INST_0_64470 : AND3
      port map(A => HIEFFPLA_NET_0_73588, B => 
        HIEFFPLA_NET_0_73587, C => HIEFFPLA_NET_0_73599, Y => 
        HIEFFPLA_NET_0_73620);
    
    HIEFFPLA_INST_0_60940 : OA1C
      port map(A => HIEFFPLA_NET_0_74338, B => 
        \General_Controller_0/flight_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_74336, Y => HIEFFPLA_NET_0_74315);
    
    \Communications_0/UART_1/rx_byte[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75378, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75496, Q => 
        \Communications_0/UART_1/rx_byte[0]_net_1\);
    
    HIEFFPLA_INST_0_70385 : AND3
      port map(A => \Timekeeper_0_microseconds[0]\, B => 
        \Timekeeper_0_microseconds[1]\, C => 
        \Timekeeper_0_microseconds[2]\, Y => HIEFFPLA_NET_0_72154);
    
    HIEFFPLA_INST_0_61821 : XA1B
      port map(A => HIEFFPLA_NET_0_73538, B => 
        \General_Controller_0/sweep_table_write_wait[1]_net_1\, C
         => HIEFFPLA_NET_0_73806, Y => HIEFFPLA_NET_0_74122);
    
    HIEFFPLA_INST_0_70300 : AND3A
      port map(A => HIEFFPLA_NET_0_72199, B => 
        HIEFFPLA_NET_0_72285, C => HIEFFPLA_NET_0_72268, Y => 
        HIEFFPLA_NET_0_72179);
    
    HIEFFPLA_INST_0_63004 : OR3B
      port map(A => HIEFFPLA_NET_0_74094, B => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, C => 
        HIEFFPLA_NET_0_73889, Y => HIEFFPLA_NET_0_73849);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72338, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\);
    
    \General_Controller_0/uc_tx_state[2]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73571, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[2]_net_1\);
    
    HIEFFPLA_INST_0_68535 : AND2
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[5]_net_1\, B => 
        GYRO_SCL_c, Y => HIEFFPLA_NET_0_72624);
    
    HIEFFPLA_INST_0_64572 : AND3C
      port map(A => HIEFFPLA_NET_0_73598, B => 
        \General_Controller_0/uc_tx_state[12]_net_1\, C => 
        \General_Controller_0/uc_tx_state[14]_net_1\, Y => 
        HIEFFPLA_NET_0_73599);
    
    HIEFFPLA_INST_0_59798 : NOR3B
      port map(A => HIEFFPLA_NET_0_74433, B => 
        HIEFFPLA_NET_0_74363, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74507);
    
    \Communications_0/UART_0/rx_byte[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75380, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75609, Q => 
        \Communications_0/UART_0/rx_byte[3]_net_1\);
    
    HIEFFPLA_INST_0_60003 : MX2
      port map(A => HIEFFPLA_NET_0_74342, B => 
        HIEFFPLA_NET_0_74402, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74475);
    
    HIEFFPLA_INST_0_67271 : AND3
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        B => HIEFFPLA_NET_0_72743, C => 
        \Sensors_0/Accelerometer_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72922);
    
    \General_Controller_0/uc_send[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73764, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73601, Q => 
        \General_Controller_0_uc_send[5]\);
    
    \General_Controller_0/sweep_table_points[6]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[6]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73981, Q => 
        \General_Controller_0/sweep_table_points[6]_net_1\);
    
    HIEFFPLA_INST_0_65067 : NAND3C
      port map(A => CLKINT_1_Y, B => HIEFFPLA_NET_0_73479, C => 
        \Pressure_Signal_Debounce_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73477);
    
    HIEFFPLA_INST_0_59692 : NOR2A
      port map(A => HIEFFPLA_NET_0_74443, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74521);
    
    HIEFFPLA_INST_0_59470 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[56]\, B => 
        \Data_Hub_Packets_0_status_packet[60]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74550);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[0]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75268, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[0]\\\\\);
    
    HIEFFPLA_INST_0_58909 : NOR3B
      port map(A => HIEFFPLA_NET_0_74371, B => 
        HIEFFPLA_NET_0_74552, C => HIEFFPLA_NET_0_74372, Y => 
        HIEFFPLA_NET_0_74661);
    
    HIEFFPLA_INST_0_59415 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[51]\, B => 
        \Data_Hub_Packets_0_status_packet[55]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74557);
    
    HIEFFPLA_INST_0_61781 : AX1C
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[1]_net_1\, B
         => \General_Controller_0/sweep_table_sweep_cnt[0]_net_1\, 
        C => 
        \General_Controller_0/sweep_table_sweep_cnt[2]_net_1\, Y
         => HIEFFPLA_NET_0_74136);
    
    \Communications_0/UART_1/tx_byte[7]\ : DFN1E1
      port map(D => \General_Controller_0_uc_send[7]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_75385, Q => 
        \Communications_0/UART_1/tx_byte[7]_net_1\);
    
    HIEFFPLA_INST_0_70688 : AX1C
      port map(A => HIEFFPLA_NET_0_72037, B => 
        \Timing_0/s_time[8]_net_1\, C => \s_clks_net_0[24]\, Y
         => HIEFFPLA_NET_0_72043);
    
    \General_Controller_0/constant_bias_probe_id[5]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73923, Q => 
        \General_Controller_0/un10_uc_tx_rdy_i[5]\);
    
    HIEFFPLA_INST_0_65708 : AX1C
      port map(A => \Science_0/ADC_READ_0/cnt4up[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt4up[0]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt4up[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73303);
    
    HIEFFPLA_INST_0_63206 : AND2B
      port map(A => HIEFFPLA_NET_0_73785, B => 
        \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73807);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[4]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72279, Q => 
        \Sensors_0_pressure_temp_raw[4]\);
    
    HIEFFPLA_INST_0_57438 : AND2
      port map(A => \Sensors_0_acc_z[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        Y => HIEFFPLA_NET_0_75046);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[15]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[15]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[15]\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73036, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_58310 : AO1
      port map(A => \Sensors_0_mag_y[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75096, Y => HIEFFPLA_NET_0_74805);
    
    \General_Controller_0/sweep_table_samples_per_step[12]\ : 
        DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[12]_net_1\);
    
    HIEFFPLA_INST_0_70494 : AX1C
      port map(A => \Timekeeper_0_milliseconds[13]\, B => 
        HIEFFPLA_NET_0_72127, C => 
        \Timekeeper_0_milliseconds[14]\, Y => 
        HIEFFPLA_NET_0_72111);
    
    HIEFFPLA_INST_0_67604 : AND3C
      port map(A => HIEFFPLA_NET_0_72929, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        C => HIEFFPLA_NET_0_72935, Y => HIEFFPLA_NET_0_72844);
    
    HIEFFPLA_INST_0_61301 : AND2A
      port map(A => HIEFFPLA_NET_0_74217, B => 
        HIEFFPLA_NET_0_74213, Y => HIEFFPLA_NET_0_74223);
    
    HIEFFPLA_INST_0_68309 : MX2
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[1]_net_1\, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_num_bytes[1]\, S
         => \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_72684);
    
    \Sensors_0/Gyro_0/I2C_Master_0/state[5]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72608, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[5]_net_1\);
    
    HIEFFPLA_INST_0_69562 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[3]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[2]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72364);
    
    HIEFFPLA_INST_0_68045 : MX2
      port map(A => HIEFFPLA_NET_0_72742, B => 
        HIEFFPLA_NET_0_72810, S => HIEFFPLA_NET_0_72878, Y => 
        HIEFFPLA_NET_0_72746);
    
    HIEFFPLA_INST_0_67265 : NOR3B
      port map(A => HIEFFPLA_NET_0_72760, B => 
        HIEFFPLA_NET_0_72885, C => HIEFFPLA_NET_0_72717, Y => 
        HIEFFPLA_NET_0_72923);
    
    HIEFFPLA_INST_0_57681 : AO1B
      port map(A => \Sensors_0_pressure_raw[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74971, Y => HIEFFPLA_NET_0_74972);
    
    HIEFFPLA_INST_0_68026 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72750);
    
    HIEFFPLA_INST_0_62646 : OR2A
      port map(A => HIEFFPLA_NET_0_74039, B => 
        HIEFFPLA_NET_0_73952, Y => HIEFFPLA_NET_0_73938);
    
    HIEFFPLA_INST_0_64267 : MX2
      port map(A => HIEFFPLA_NET_0_73739, B => 
        HIEFFPLA_NET_0_73731, S => HIEFFPLA_NET_0_73588, Y => 
        HIEFFPLA_NET_0_73643);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[0]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72767, Q => 
        \Sensors_0_acc_y[0]\);
    
    \Science_0/ADC_READ_0/chan7_data[2]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[8]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[2]\);
    
    HIEFFPLA_INST_0_66407 : XA1C
      port map(A => HIEFFPLA_NET_0_73131, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[3]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_73127);
    
    HIEFFPLA_INST_0_64933 : MX2C
      port map(A => HIEFFPLA_NET_0_73508, B => 
        HIEFFPLA_NET_0_73518, S => 
        \I2C_PassThrough_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73509);
    
    HIEFFPLA_INST_0_65565 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt3dn[5]_net_1\, B => 
        HIEFFPLA_NET_0_73351, C => HIEFFPLA_NET_0_73349, Y => 
        HIEFFPLA_NET_0_73342);
    
    HIEFFPLA_INST_0_57444 : AOI1
      port map(A => \Science_0_exp_packet_0[26]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_75043, Y => HIEFFPLA_NET_0_75044);
    
    HIEFFPLA_INST_0_63376 : MX2
      port map(A => HIEFFPLA_NET_0_73761, B => 
        HIEFFPLA_NET_0_73697, S => HIEFFPLA_NET_0_73608, Y => 
        HIEFFPLA_NET_0_73769);
    
    HIEFFPLA_INST_0_54929 : AND2
      port map(A => TOP_UART_RX_c, B => EMU_RX_c, Y => 
        HIEFFPLA_NET_0_75638);
    
    HIEFFPLA_INST_0_71207 : AOI1B
      port map(A => HIEFFPLA_NET_0_75478, B => 
        HIEFFPLA_NET_0_75479, C => 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\, Y => 
        HIEFFPLA_NET_0_71974);
    
    HIEFFPLA_INST_0_60885 : NAND3C
      port map(A => \General_Controller_0/command[0]_net_1\, B
         => HIEFFPLA_NET_0_74329, C => HIEFFPLA_NET_0_74335, Y
         => HIEFFPLA_NET_0_74330);
    
    HIEFFPLA_INST_0_59959 : NOR3B
      port map(A => HIEFFPLA_NET_0_74556, B => 
        HIEFFPLA_NET_0_74432, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74482);
    
    \General_Controller_0/uc_rx_state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74065, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_state[0]_net_1\);
    
    HIEFFPLA_INST_0_69295 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72426);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[6]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_75247, CLK => CLKINT_0_Y_0, E
         => CLKINT_1_Y, Q => 
        \Data_Saving_0/Interrupt_Generator_0/counter[6]_net_1\);
    
    \Science_0/DAC_SET_0/vector[14]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73199, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[14]_net_1\);
    
    HIEFFPLA_INST_0_55023 : AND3
      port map(A => HIEFFPLA_NET_0_75593, B => 
        HIEFFPLA_NET_0_75591, C => HIEFFPLA_NET_0_75603, Y => 
        HIEFFPLA_NET_0_75612);
    
    HIEFFPLA_INST_0_67359 : NOR3B
      port map(A => HIEFFPLA_NET_0_72888, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, C
         => HIEFFPLA_NET_0_72791, Y => HIEFFPLA_NET_0_72899);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[8]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72283, Q => 
        \Sensors_0_pressure_temp_raw[8]\);
    
    HIEFFPLA_INST_0_66485 : MIN3X
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73109);
    
    HIEFFPLA_INST_0_65331 : XA1B
      port map(A => \Science_0/ADC_READ_0/cnt1dn[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt1dn[0]_net_1\, C => 
        HIEFFPLA_NET_0_73244, Y => HIEFFPLA_NET_0_73407);
    
    HIEFFPLA_INST_0_69359 : MX2
      port map(A => HIEFFPLA_NET_0_72404, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_num_bytes[0]\, 
        S => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72408);
    
    HIEFFPLA_INST_0_56080 : AND3
      port map(A => HIEFFPLA_NET_0_75351, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\, C
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, 
        Y => HIEFFPLA_NET_0_75352);
    
    HIEFFPLA_INST_0_56539 : XOR2
      port map(A => HIEFFPLA_NET_0_75255, B => 
        \Data_Saving_0/Interrupt_Generator_0/counter[7]_net_1\, Y
         => HIEFFPLA_NET_0_75246);
    
    HIEFFPLA_INST_0_68824 : OR2A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, B
         => CLKINT_1_Y, Y => HIEFFPLA_NET_0_72548);
    
    HIEFFPLA_INST_0_62991 : NAND3C
      port map(A => HIEFFPLA_NET_0_73829, B => 
        HIEFFPLA_NET_0_73826, C => HIEFFPLA_NET_0_74008, Y => 
        HIEFFPLA_NET_0_73851);
    
    HIEFFPLA_INST_0_69114 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[2]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[1]_net_1\, 
        C => HIEFFPLA_NET_0_72557, Y => HIEFFPLA_NET_0_72468);
    
    HIEFFPLA_INST_0_64031 : MX2
      port map(A => HIEFFPLA_NET_0_73641, B => 
        HIEFFPLA_NET_0_73633, S => HIEFFPLA_NET_0_73585, Y => 
        HIEFFPLA_NET_0_73678);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/data_out[6]\ : 
        DFN0E1C1
      port map(D => PRESSURE_SDA_in, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72396, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[6]\);
    
    HIEFFPLA_INST_0_62723 : AND3C
      port map(A => HIEFFPLA_NET_0_73788, B => 
        HIEFFPLA_NET_0_73804, C => 
        \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73921);
    
    HIEFFPLA_INST_0_58903 : AND2B
      port map(A => HIEFFPLA_NET_0_74636, B => 
        \GS_Readout_0/state[0]_net_1\, Y => HIEFFPLA_NET_0_74662);
    
    HIEFFPLA_INST_0_66161 : MX2B
      port map(A => \Science_0/DAC_SET_0/vector[2]_net_1\, B => 
        \Science_0/DAC_SET_0/ADR[1]_net_1\, S => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73193);
    
    HIEFFPLA_INST_0_57615 : AO1B
      port map(A => \Sensors_0_gyro_x[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74991, Y => HIEFFPLA_NET_0_74992);
    
    HIEFFPLA_INST_0_55603 : AND2B
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[25]_net_1\, B => 
        \Communications_0/UART_1/rx_clk_count[26]_net_1\, Y => 
        HIEFFPLA_NET_0_75468);
    
    HIEFFPLA_INST_0_62091 : AO1A
      port map(A => HIEFFPLA_NET_0_73875, B => 
        \General_Controller_0/uc_rx_prev_state[4]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74054);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[11]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72484, Q => 
        \Sensors_0_gyro_y[11]\);
    
    HIEFFPLA_INST_0_62012 : NOR2A
      port map(A => \General_Controller_0/uc_rx_byte[5]_net_1\, B
         => \General_Controller_0/uc_rx_byte[6]_net_1\, Y => 
        HIEFFPLA_NET_0_74074);
    
    HIEFFPLA_INST_0_61109 : AO1
      port map(A => HIEFFPLA_NET_0_74282, B => 
        \Timekeeper_0_milliseconds[3]\, C => 
        \Timekeeper_0_milliseconds[4]\, Y => HIEFFPLA_NET_0_74274);
    
    \Communications_0/FFU_Command_Checker_0/command_out[2]\ : 
        DFN1E1C1
      port map(D => \Communications_0/UART_0_recv[2]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75625, Q => \Communications_0_ext_recv[2]\);
    
    HIEFFPLA_INST_0_62833 : AND2
      port map(A => \General_Controller_0/uc_rx_state[4]_net_1\, 
        B => \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73888);
    
    HIEFFPLA_INST_0_58485 : OA1A
      port map(A => General_Controller_0_en_data_saving, B => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, C => 
        HIEFFPLA_NET_0_74752, Y => HIEFFPLA_NET_0_74753);
    
    \General_Controller_0/st_raddr[2]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[2]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73979, Q => 
        \General_Controller_0_st_raddr_1[2]\);
    
    HIEFFPLA_INST_0_67684 : NOR3B
      port map(A => HIEFFPLA_NET_0_72743, B => 
        HIEFFPLA_NET_0_72820, C => HIEFFPLA_NET_0_72792, Y => 
        HIEFFPLA_NET_0_72824);
    
    HIEFFPLA_INST_0_55595 : NOR3B
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[28]_net_1\, B => 
        \Communications_0/UART_1/rx_clk_count[27]_net_1\, C => 
        HIEFFPLA_NET_0_75467, Y => HIEFFPLA_NET_0_75470);
    
    HIEFFPLA_INST_0_68793 : AND2B
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0_write_done\, B
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        Y => HIEFFPLA_NET_0_72560);
    
    HIEFFPLA_INST_0_70559 : AND2B
      port map(A => \Timing_0/m_count[0]_net_1\, B => 
        HIEFFPLA_NET_0_72083, Y => HIEFFPLA_NET_0_72080);
    
    HIEFFPLA_INST_0_65412 : OR3A
      port map(A => \Science_0/ADC_READ_0/cnt2dn[3]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2dn[5]_net_1\, C => 
        HIEFFPLA_NET_0_73378, Y => HIEFFPLA_NET_0_73383);
    
    \General_Controller_0/constant_bias_voltage_1[11]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[11]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/packet_select[5]\ : DFN0E0C1
      port map(D => 
        \Data_Saving_0/Packet_Saver_0/ch_0_flag_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\);
    
    \ACLK_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => ACLK_c, E => \VCC\, DOUT => 
        \ACLK_pad/U0/NET1\, EOUT => \ACLK_pad/U0/NET2\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/data_out_1[0]\ : 
        DFN1E1
      port map(D => HIEFFPLA_NET_0_73007, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72795, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[0]\);
    
    HIEFFPLA_INST_0_88376 : XOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[7]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[8]\\\\\, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[10]\\\\\, Y
         => HIEFFPLA_NET_0_88382);
    
    HIEFFPLA_INST_0_66785 : NOR3A
      port map(A => HIEFFPLA_NET_0_73034, B => 
        HIEFFPLA_NET_0_73020, C => HIEFFPLA_NET_0_73023, Y => 
        HIEFFPLA_NET_0_73035);
    
    HIEFFPLA_INST_0_71068 : MX2
      port map(A => \GS_Readout_0/state[4]_net_1\, B => 
        \GS_Readout_0/state[3]_net_1\, S => HIEFFPLA_NET_0_74382, 
        Y => HIEFFPLA_NET_0_71982);
    
    HIEFFPLA_INST_0_57953 : AO1
      port map(A => \Science_0_exp_packet_0[70]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75163, Y => HIEFFPLA_NET_0_74895);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72870, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\);
    
    HIEFFPLA_INST_0_62966 : NOR2A
      port map(A => \General_Controller_0/uc_rx_state[3]_net_1\, 
        B => HIEFFPLA_NET_0_73855, Y => HIEFFPLA_NET_0_73856);
    
    HIEFFPLA_INST_0_69631 : AO1
      port map(A => HIEFFPLA_NET_0_72349, B => 
        HIEFFPLA_NET_0_72390, C => HIEFFPLA_NET_0_72339, Y => 
        HIEFFPLA_NET_0_72340);
    
    HIEFFPLA_INST_0_66272 : NAND3
      port map(A => HIEFFPLA_NET_0_73159, B => 
        HIEFFPLA_NET_0_73161, C => HIEFFPLA_NET_0_73157, Y => 
        HIEFFPLA_NET_0_73160);
    
    HIEFFPLA_INST_0_60420 : MX2
      port map(A => \Science_0_chan7_data[8]\, B => 
        \Science_0_chan6_data[0]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74418);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/s_ack_error\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72347, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72385, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_s_ack_error\);
    
    HIEFFPLA_INST_0_56281 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[10]\\\\\, B
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[9]\\\\\, Y
         => HIEFFPLA_NET_0_75320);
    
    \Science_0/ADC_READ_0/exp_packet_1[65]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[9]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[65]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/data_out_1[6]\ : 
        DFN1E1
      port map(D => HIEFFPLA_NET_0_73002, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72795, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[6]\);
    
    HIEFFPLA_INST_0_61191 : AND2
      port map(A => 
        \General_Controller_0/state_seconds[17]_net_1\, B => 
        \General_Controller_0/state_seconds[16]_net_1\, Y => 
        HIEFFPLA_NET_0_74254);
    
    HIEFFPLA_INST_0_68201 : NOR2A
      port map(A => \Sensors_0/Accelerometer_0/state[8]\, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72708);
    
    HIEFFPLA_INST_0_66950 : AND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_72793, Y => HIEFFPLA_NET_0_72998);
    
    HIEFFPLA_INST_0_55348 : OR2A
      port map(A => HIEFFPLA_NET_0_75534, B => 
        \Communications_0/UART_0/tx_clk_count_i_0[6]\, Y => 
        HIEFFPLA_NET_0_75535);
    
    HIEFFPLA_INST_0_61265 : AX1
      port map(A => HIEFFPLA_NET_0_74244, B => 
        \General_Controller_0/state_seconds[14]_net_1\, C => 
        \General_Controller_0/state_seconds[15]_net_1\, Y => 
        HIEFFPLA_NET_0_74233);
    
    HIEFFPLA_INST_0_55829 : NAND3C
      port map(A => HIEFFPLA_NET_0_75386, B => 
        HIEFFPLA_NET_0_75417, C => 
        \Communications_0/UART_1/tx_clk_count_i_0[2]\, Y => 
        HIEFFPLA_NET_0_75418);
    
    HIEFFPLA_INST_0_70241 : OR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[4]_net_1\, 
        C => HIEFFPLA_NET_0_72240, Y => HIEFFPLA_NET_0_72188);
    
    HIEFFPLA_INST_0_61977 : AND2B
      port map(A => \General_Controller_0/uc_rx_byte[1]_net_1\, B
         => \General_Controller_0/uc_rx_byte[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74085);
    
    HIEFFPLA_INST_0_60549 : NOR2A
      port map(A => HIEFFPLA_NET_0_74556, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74397);
    
    \GS_Readout_0/state[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74607, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/state[3]_net_1\);
    
    \SweepTable_0/SweepTable_R0C0\ : RAM512X18
      port map(RADDR8 => AFLSDF_GND, RADDR7 => 
        \TableSelect_0_RADDR[7]\, RADDR6 => 
        \TableSelect_0_RADDR[6]\, RADDR5 => 
        \TableSelect_0_RADDR[5]\, RADDR4 => 
        \TableSelect_0_RADDR[4]\, RADDR3 => 
        \TableSelect_0_RADDR[3]\, RADDR2 => 
        \TableSelect_0_RADDR[2]\, RADDR1 => 
        \TableSelect_0_RADDR[1]\, RADDR0 => 
        \TableSelect_0_RADDR[0]\, WADDR8 => AFLSDF_GND, WADDR7
         => \General_Controller_0_st_waddr[7]\, WADDR6 => 
        \General_Controller_0_st_waddr[6]\, WADDR5 => 
        \General_Controller_0_st_waddr[5]\, WADDR4 => 
        \General_Controller_0_st_waddr[4]\, WADDR3 => 
        \General_Controller_0_st_waddr[3]\, WADDR2 => 
        \General_Controller_0_st_waddr[2]\, WADDR1 => 
        \General_Controller_0_st_waddr[1]\, WADDR0 => 
        \General_Controller_0_st_waddr[0]\, WD17 => \GND\, WD16
         => \General_Controller_0_st_wdata[15]\, WD15 => 
        \General_Controller_0_st_wdata[14]\, WD14 => 
        \General_Controller_0_st_wdata[13]\, WD13 => 
        \General_Controller_0_st_wdata[12]\, WD12 => 
        \General_Controller_0_st_wdata[11]\, WD11 => 
        \General_Controller_0_st_wdata[10]\, WD10 => 
        \General_Controller_0_st_wdata[9]\, WD9 => 
        \General_Controller_0_st_wdata[8]\, WD8 => \GND\, WD7 => 
        \General_Controller_0_st_wdata[7]\, WD6 => 
        \General_Controller_0_st_wdata[6]\, WD5 => 
        \General_Controller_0_st_wdata[5]\, WD4 => 
        \General_Controller_0_st_wdata[4]\, WD3 => 
        \General_Controller_0_st_wdata[3]\, WD2 => 
        \General_Controller_0_st_wdata[2]\, WD1 => 
        \General_Controller_0_st_wdata[1]\, WD0 => 
        \General_Controller_0_st_wdata[0]\, RW0 => \GND\, RW1 => 
        \VCC\, WW0 => \GND\, WW1 => \VCC\, PIPE => \VCC\, REN => 
        \AFLSDF_INV_4\, WEN => \SweepTable_0.WEAP\, RCLK => 
        CLKINT_0_Y_0, WCLK => CLKINT_0_Y_0, RESET => 
        \AFLSDF_INV_5\, RD17 => OPEN, RD16 => 
        \SweepTable_0_RD[15]\, RD15 => \SweepTable_0_RD[14]\, 
        RD14 => \SweepTable_0_RD[13]\, RD13 => 
        \SweepTable_0_RD[12]\, RD12 => \SweepTable_0_RD[11]\, 
        RD11 => \SweepTable_0_RD[10]\, RD10 => 
        \SweepTable_0_RD[9]\, RD9 => \SweepTable_0_RD[8]\, RD8
         => OPEN, RD7 => \SweepTable_0_RD[7]\, RD6 => 
        \SweepTable_0_RD[6]\, RD5 => \SweepTable_0_RD[5]\, RD4
         => \SweepTable_0_RD[4]\, RD3 => \SweepTable_0_RD[3]\, 
        RD2 => \SweepTable_0_RD[2]\, RD1 => \SweepTable_0_RD[1]\, 
        RD0 => \SweepTable_0_RD[0]\);
    
    HIEFFPLA_INST_0_66439 : NAND3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        C => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73121);
    
    HIEFFPLA_INST_0_60963 : AO1A
      port map(A => HIEFFPLA_NET_0_74313, B => 
        HIEFFPLA_NET_0_74308, C => HIEFFPLA_NET_0_74307, Y => 
        HIEFFPLA_NET_0_74309);
    
    HIEFFPLA_INST_0_55013 : XO1
      port map(A => \General_Controller_0_unit_id[2]\, B => 
        \Communications_0/UART_0_recv[2]\, C => 
        HIEFFPLA_NET_0_75615, Y => HIEFFPLA_NET_0_75616);
    
    HIEFFPLA_INST_0_70507 : AX1C
      port map(A => \Timekeeper_0_milliseconds[19]\, B => 
        HIEFFPLA_NET_0_72123, C => 
        \Timekeeper_0_milliseconds[20]\, Y => 
        HIEFFPLA_NET_0_72104);
    
    \Data_Saving_0/Packet_Saver_0/data_out[12]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75233, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[12]\);
    
    HIEFFPLA_INST_0_69593 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[5]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72355);
    
    HIEFFPLA_INST_0_68975 : AOI1
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, B
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        C => \Sensors_0/Gyro_0/I2C_Master_0_s_ack_error\, Y => 
        HIEFFPLA_NET_0_72509);
    
    HIEFFPLA_INST_0_56401 : XOR2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[6]\\\\\, B
         => HIEFFPLA_NET_0_75348, Y => HIEFFPLA_NET_0_75288);
    
    HIEFFPLA_INST_0_59807 : NOR3A
      port map(A => \GS_Readout_0/subState[2]_net_1\, B => 
        \GS_Readout_0/subState[0]_net_1\, C => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74505);
    
    HIEFFPLA_INST_0_57900 : AOI1
      port map(A => \Sensors_0_acc_time[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74910, Y => HIEFFPLA_NET_0_74911);
    
    HIEFFPLA_INST_0_64892 : XA1
      port map(A => HIEFFPLA_NET_0_73503, B => 
        \I2C_PassThrough_0/cnt[4]_net_1\, C => 
        HIEFFPLA_NET_0_73515, Y => HIEFFPLA_NET_0_73516);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[11]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[11]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[11]\);
    
    HIEFFPLA_INST_0_68254 : XAI1A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, B => 
        HIEFFPLA_NET_0_72574, C => HIEFFPLA_NET_0_72622, Y => 
        HIEFFPLA_NET_0_72696);
    
    HIEFFPLA_INST_0_69791 : AO1E
      port map(A => HIEFFPLA_NET_0_72308, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[0]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72302);
    
    HIEFFPLA_INST_0_63075 : MX2
      port map(A => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        B => \General_Controller_0/uc_rx_byte[3]_net_1\, S => 
        \General_Controller_0/uc_rx_byte[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73835);
    
    HIEFFPLA_INST_0_62806 : NAND3C
      port map(A => HIEFFPLA_NET_0_73854, B => 
        HIEFFPLA_NET_0_73960, C => HIEFFPLA_NET_0_73892, Y => 
        HIEFFPLA_NET_0_73898);
    
    HIEFFPLA_INST_0_57192 : AO1
      port map(A => \Sensors_0_mag_time[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75093, Y => HIEFFPLA_NET_0_75134);
    
    HIEFFPLA_INST_0_68537 : NAND3C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_72623);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[12]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72490, Q => 
        \ch3_data_net_0[8]\);
    
    HIEFFPLA_INST_0_69175 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        B => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, 
        C => \Sensors_0/Gyro_0/I2C_Master_0_write_done\, Y => 
        HIEFFPLA_NET_0_72455);
    
    HIEFFPLA_INST_0_66506 : AOI1
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_73106);
    
    HIEFFPLA_INST_0_55836 : AND3
      port map(A => \Communications_0/UART_1/tx_clk_count_i_0[5]\, 
        B => \Communications_0/UART_1/tx_clk_count_i_0[7]\, C => 
        \Communications_0/UART_1/tx_clk_count_i_0[6]\, Y => 
        HIEFFPLA_NET_0_75415);
    
    \General_Controller_0/sweep_table_samples_per_point[15]\ : 
        DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[15]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[9]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72800, Q => 
        \Sensors_0_acc_x[9]\);
    
    \Science_0/ADC_READ_0/chan6_data[9]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[9]\);
    
    \Science_0/ADC_READ_0/chan0_data[9]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[9]\);
    
    HIEFFPLA_INST_0_64357 : MX2
      port map(A => HIEFFPLA_NET_0_73722, B => 
        HIEFFPLA_NET_0_73714, S => HIEFFPLA_NET_0_73619, Y => 
        HIEFFPLA_NET_0_73634);
    
    HIEFFPLA_INST_0_62265 : AO1
      port map(A => HIEFFPLA_NET_0_74153, B => 
        HIEFFPLA_NET_0_73972, C => HIEFFPLA_NET_0_74127, Y => 
        HIEFFPLA_NET_0_74017);
    
    HIEFFPLA_INST_0_59812 : MX2
      port map(A => \ch3_data_net_0[2]\, B => \ch3_data_net_0[6]\, 
        S => \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74504);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72534, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[5]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72777, Q => 
        \Sensors_0_acc_y[5]\);
    
    HIEFFPLA_INST_0_67646 : NOR3B
      port map(A => HIEFFPLA_NET_0_72743, B => 
        HIEFFPLA_NET_0_72882, C => HIEFFPLA_NET_0_72792, Y => 
        HIEFFPLA_NET_0_72834);
    
    \Timing_0/m_count[4]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72076, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_count[4]_net_1\);
    
    HIEFFPLA_INST_0_57038 : MX2
      port map(A => HIEFFPLA_NET_0_74954, B => 
        HIEFFPLA_NET_0_74768, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75178);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[7]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72777, Q => 
        \Sensors_0_acc_y[7]\);
    
    HIEFFPLA_INST_0_62344 : AO1A
      port map(A => HIEFFPLA_NET_0_73788, B => 
        HIEFFPLA_NET_0_73913, C => HIEFFPLA_NET_0_74004, Y => 
        HIEFFPLA_NET_0_74001);
    
    HIEFFPLA_INST_0_71061 : AND3C
      port map(A => HIEFFPLA_NET_0_71984, B => 
        \General_Controller_0/state_seconds[7]_net_1\, C => 
        \General_Controller_0/state_seconds[6]_net_1\, Y => 
        HIEFFPLA_NET_0_74252);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[6]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72276, Q => \Sensors_0_pressure_raw[6]\);
    
    HIEFFPLA_INST_0_67981 : AND3
      port map(A => \Sensors_0/Accelerometer_0/state[8]\, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72762);
    
    HIEFFPLA_INST_0_65570 : XA1
      port map(A => HIEFFPLA_NET_0_73358, B => 
        \Science_0/ADC_READ_0/cnt3dn[6]_net_1\, C => 
        HIEFFPLA_NET_0_73349, Y => HIEFFPLA_NET_0_73341);
    
    HIEFFPLA_INST_0_70794 : AO1A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, B
         => HIEFFPLA_NET_0_72010, C => HIEFFPLA_NET_0_72478, Y
         => HIEFFPLA_NET_0_72432);
    
    HIEFFPLA_INST_0_65478 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt2up[0]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2up[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt2up[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73367);
    
    \Science_0/DAC_SET_0/vector[9]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73187, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[9]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/data_out_1[3]\ : 
        DFN1E1
      port map(D => HIEFFPLA_NET_0_73005, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72795, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[3]\);
    
    HIEFFPLA_INST_0_55482 : AND2B
      port map(A => \Communications_0/UART_0/tx_state[0]_net_1\, 
        B => \Communications_0/UART_0/tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75501);
    
    HIEFFPLA_INST_0_69245 : AND3
      port map(A => HIEFFPLA_NET_0_72438, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, C
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        Y => HIEFFPLA_NET_0_72440);
    
    HIEFFPLA_INST_0_60949 : NAND2
      port map(A => \Timekeeper_0_milliseconds[6]\, B => 
        \Timekeeper_0_milliseconds[5]\, Y => HIEFFPLA_NET_0_74313);
    
    HIEFFPLA_INST_0_57430 : AND2
      port map(A => \Sensors_0_gyro_temp[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75048);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_READ_RESET_P\ : DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_2_Q\, CLK
         => CLKINT_2_Y, CLR => \AFLSDF_INV_31\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\);
    
    HIEFFPLA_INST_0_55131 : AND2B
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[23]_net_1\, B => 
        \Communications_0/UART_0/rx_clk_count[24]_net_1\, Y => 
        HIEFFPLA_NET_0_75580);
    
    HIEFFPLA_INST_0_66813 : AO1A
      port map(A => HIEFFPLA_NET_0_73098, B => 
        HIEFFPLA_NET_0_73026, C => HIEFFPLA_NET_0_73022, Y => 
        HIEFFPLA_NET_0_73029);
    
    HIEFFPLA_INST_0_67081 : AO1A
      port map(A => HIEFFPLA_NET_0_72752, B => 
        HIEFFPLA_NET_0_72925, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/isSetup_net_1\, 
        Y => HIEFFPLA_NET_0_72969);
    
    \General_Controller_0/constant_bias_voltage_1[13]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[13]_net_1\);
    
    HIEFFPLA_INST_0_62077 : AO1D
      port map(A => HIEFFPLA_NET_0_73862, B => 
        \General_Controller_0/uc_rx_state_0[1]_net_1\, C => 
        HIEFFPLA_NET_0_74052, Y => HIEFFPLA_NET_0_74057);
    
    HIEFFPLA_INST_0_57937 : AO1B
      port map(A => \Sensors_0_gyro_time[13]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74899, Y => HIEFFPLA_NET_0_74900);
    
    HIEFFPLA_INST_0_67006 : AOI1D
      port map(A => HIEFFPLA_NET_0_72890, B => 
        HIEFFPLA_NET_0_72913, C => HIEFFPLA_NET_0_72735, Y => 
        HIEFFPLA_NET_0_72986);
    
    \Data_Saving_0/Interrupt_Generator_0/counter[3]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_75250, CLK => CLKINT_0_Y_0, E
         => CLKINT_1_Y, Q => 
        \Data_Saving_0/Interrupt_Generator_0/counter[3]_net_1\);
    
    HIEFFPLA_INST_0_57877 : AO1B
      port map(A => \Sensors_0_mag_time[23]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74917, Y => HIEFFPLA_NET_0_74918);
    
    \Data_Saving_0/Packet_Saver_0/pressure_flag\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_74765, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => 
        General_Controller_0_en_data_saving, Q => 
        \Data_Saving_0/Packet_Saver_0/pressure_flag_net_1\);
    
    HIEFFPLA_INST_0_59013 : AO1C
      port map(A => HIEFFPLA_NET_0_74360, B => 
        HIEFFPLA_NET_0_74368, C => \GS_Readout_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_74637);
    
    HIEFFPLA_INST_0_69024 : AO1E
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        B => HIEFFPLA_NET_0_72493, C => HIEFFPLA_NET_0_72540, Y
         => HIEFFPLA_NET_0_72494);
    
    \GS_Readout_0/prevState[3]\ : DFN1E0C1
      port map(D => \GS_Readout_0/state[3]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \GS_Readout_0/state[6]_net_1\, Q => 
        \GS_Readout_0/prevState[3]_net_1\);
    
    \General_Controller_0/st_waddr[7]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_waddr[7]\);
    
    AFLSDF_INV_12 : INV
      port map(A => CLKINT_1_Y, Y => \AFLSDF_INV_12\);
    
    HIEFFPLA_INST_0_62903 : OA1A
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73870);
    
    HIEFFPLA_INST_0_61306 : XA1C
      port map(A => HIEFFPLA_NET_0_74248, B => 
        \General_Controller_0/state_seconds[5]_net_1\, C => 
        HIEFFPLA_NET_0_74217, Y => HIEFFPLA_NET_0_74222);
    
    \General_Controller_0/status_bits_1[49]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74197, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[49]\);
    
    \General_Controller_0/command[7]\ : DFN1E1
      port map(D => \Communications_0_ext_recv[7]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74300, Q => 
        \General_Controller_0/command[7]_net_1\);
    
    HIEFFPLA_INST_0_68990 : OR2A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        B => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72505);
    
    HIEFFPLA_INST_0_61761 : XOR2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[0]_net_1\, B
         => HIEFFPLA_NET_0_73927, Y => HIEFFPLA_NET_0_74144);
    
    HIEFFPLA_INST_0_68772 : MX2B
      port map(A => HIEFFPLA_NET_0_72488, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, S
         => HIEFFPLA_NET_0_72539, Y => HIEFFPLA_NET_0_72565);
    
    \Science_0/DAC_SET_0/vector[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73192, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[4]_net_1\);
    
    \Timekeeper_0/microseconds[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72151, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timekeeper_0_microseconds[0]\);
    
    HIEFFPLA_INST_0_56278 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[5]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[4]\\\\\, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[3]\\\\\, Y => 
        HIEFFPLA_NET_0_75322);
    
    HIEFFPLA_INST_0_70563 : AOI1B
      port map(A => HIEFFPLA_NET_0_72082, B => 
        HIEFFPLA_NET_0_72081, C => HIEFFPLA_NET_0_72078, Y => 
        HIEFFPLA_NET_0_72079);
    
    HIEFFPLA_INST_0_63788 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[2]_net_1\, 
        B => \General_Controller_0/sweep_table_points[2]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73711);
    
    HIEFFPLA_INST_0_57618 : AOI1
      port map(A => \Science_0_exp_packet_0[46]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74798, Y => HIEFFPLA_NET_0_74991);
    
    HIEFFPLA_INST_0_60879 : NOR3B
      port map(A => HIEFFPLA_NET_0_74331, B => 
        \General_Controller_0/command[3]_net_1\, C => 
        \General_Controller_0/ext_rx_state_i_0[1]\, Y => 
        HIEFFPLA_NET_0_74332);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[8]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72777, Q => 
        \Sensors_0_acc_y[8]\);
    
    HIEFFPLA_INST_0_69775 : AND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[6]_net_1\, 
        Y => HIEFFPLA_NET_0_72310);
    
    HIEFFPLA_INST_0_60988 : OR2A
      port map(A => HIEFFPLA_NET_0_74339, B => 
        \General_Controller_0/flight_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74303);
    
    HIEFFPLA_INST_0_58274 : AO1
      port map(A => \Sensors_0_gyro_time[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75108, Y => HIEFFPLA_NET_0_74814);
    
    HIEFFPLA_INST_0_58209 : AND2
      port map(A => \Sensors_0_pressure_temp_raw[14]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_74828);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]\ : 
        DFN1P1
      port map(D => HIEFFPLA_NET_0_72261, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\);
    
    \General_Controller_0/command[3]\ : DFN1E1
      port map(D => \Communications_0_ext_recv[3]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74300, Q => 
        \General_Controller_0/command[3]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[19]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[3]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[19]\);
    
    HIEFFPLA_INST_0_62901 : OA1C
      port map(A => HIEFFPLA_NET_0_74027, B => 
        HIEFFPLA_NET_0_73781, C => HIEFFPLA_NET_0_73946, Y => 
        HIEFFPLA_NET_0_73871);
    
    HIEFFPLA_INST_0_66692 : AO1A
      port map(A => ACCE_SDA_in, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        C => CLKINT_1_Y, Y => HIEFFPLA_NET_0_73062);
    
    HIEFFPLA_INST_0_57990 : NAND3C
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        C => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_74885);
    
    HIEFFPLA_INST_0_62563 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state[1]_net_1\, 
        B => \General_Controller_0/uc_rx_state[3]_net_1\, C => 
        HIEFFPLA_NET_0_73909, Y => HIEFFPLA_NET_0_73956);
    
    HIEFFPLA_INST_0_63308 : OR3B
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, C => 
        HIEFFPLA_NET_0_73785, Y => HIEFFPLA_NET_0_73781);
    
    HIEFFPLA_INST_0_60605 : AND3
      port map(A => HIEFFPLA_NET_0_74341, B => 
        HIEFFPLA_NET_0_74342, C => HIEFFPLA_NET_0_74546, Y => 
        HIEFFPLA_NET_0_74388);
    
    \General_Controller_0/state_seconds[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74221, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[6]_net_1\);
    
    HIEFFPLA_INST_0_65323 : AND2B
      port map(A => \Science_0/ADC_READ_0/cnt1dn[5]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt1dn[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73411);
    
    HIEFFPLA_INST_0_57863 : AO1
      port map(A => \Science_0_exp_packet_0[77]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75138, Y => HIEFFPLA_NET_0_74922);
    
    \GYRO_SDA_pad/U0/U1\ : IOBI_IB_OB_EB
      port map(D => \Sensors_0.Gyro_0.I2C_Master_0.sda_1\, E => 
        sda_cl_1_RNITJT01, YIN => \GYRO_SDA_pad/U0/NET3\, DOUT
         => \GYRO_SDA_pad/U0/NET1\, EOUT => 
        \GYRO_SDA_pad/U0/NET2\, Y => GYRO_SDA_in);
    
    HIEFFPLA_INST_0_56568 : AND2
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/old_ch_0_new_data_i_0\, B
         => Science_0_exp_new_data, Y => HIEFFPLA_NET_0_75237);
    
    \Communications_0/UART_1/tx_byte[2]\ : DFN1E1
      port map(D => \General_Controller_0_uc_send[2]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_75385, Q => 
        \Communications_0/UART_1/tx_byte[2]_net_1\);
    
    HIEFFPLA_INST_0_57647 : AO1
      port map(A => \Sensors_0_pressure_raw[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74793, Y => HIEFFPLA_NET_0_74982);
    
    \Science_0/ADC_READ_0/chan5_data[1]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[1]\);
    
    HIEFFPLA_INST_0_58874 : AOI1
      port map(A => HIEFFPLA_NET_0_74698, B => 
        HIEFFPLA_NET_0_74569, C => HIEFFPLA_NET_0_74696, Y => 
        HIEFFPLA_NET_0_74668);
    
    HIEFFPLA_INST_0_55029 : AND3
      port map(A => HIEFFPLA_NET_0_75593, B => 
        HIEFFPLA_NET_0_75591, C => HIEFFPLA_NET_0_75601, Y => 
        HIEFFPLA_NET_0_75610);
    
    \Science_0/ADC_READ_0/exp_packet_1[71]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[15]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[71]\);
    
    HIEFFPLA_INST_0_63057 : AO1A
      port map(A => HIEFFPLA_NET_0_73889, B => 
        HIEFFPLA_NET_0_73791, C => HIEFFPLA_NET_0_73833, Y => 
        HIEFFPLA_NET_0_73839);
    
    \FFU_EJECTED_pad/U0/U0\ : IOPAD_IN
      port map(PAD => FFU_EJECTED, Y => \FFU_EJECTED_pad/U0/NET1\);
    
    HIEFFPLA_INST_0_58753 : NOR3B
      port map(A => \GS_Readout_0/state[1]_net_1\, B => 
        HIEFFPLA_NET_0_74432, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74692);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72466, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[3]_net_1\);
    
    \SCIENCE_TX_pad/U0/U0\ : IOPAD_TRI
      port map(D => \SCIENCE_TX_pad/U0/NET1\, E => 
        \SCIENCE_TX_pad/U0/NET2\, PAD => SCIENCE_TX);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[6]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72808, Q => 
        \Sensors_0_mag_z[6]\);
    
    \Science_0/ADC_READ_0/chan7_data[9]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[15]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[9]\);
    
    HIEFFPLA_INST_0_65191 : AND2
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[0]_net_1\, 
        B => HIEFFPLA_NET_0_73478, Y => HIEFFPLA_NET_0_73449);
    
    HIEFFPLA_INST_0_64693 : NOR2A
      port map(A => Communications_0_uc_tx_rdy, B => 
        HIEFFPLA_NET_0_73560, Y => HIEFFPLA_NET_0_73562);
    
    HIEFFPLA_INST_0_69000 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, B
         => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        C => CLKINT_1_Y, Y => HIEFFPLA_NET_0_72502);
    
    HIEFFPLA_INST_0_61524 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[58]\, B => 
        \Timekeeper_0_milliseconds[18]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74188);
    
    HIEFFPLA_INST_0_68950 : NOR3B
      port map(A => HIEFFPLA_NET_0_72508, B => 
        HIEFFPLA_NET_0_72512, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72515);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/num_bytes_1[1]\ : 
        DFN1E1
      port map(D => HIEFFPLA_NET_0_72494, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72549, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_num_bytes[1]\);
    
    HIEFFPLA_INST_0_67210 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        B => HIEFFPLA_NET_0_72717, C => HIEFFPLA_NET_0_72744, Y
         => HIEFFPLA_NET_0_72938);
    
    HIEFFPLA_INST_0_60859 : NAND2B
      port map(A => HIEFFPLA_NET_0_74328, B => 
        HIEFFPLA_NET_0_74334, Y => HIEFFPLA_NET_0_74338);
    
    HIEFFPLA_INST_0_58706 : NOR3B
      port map(A => HIEFFPLA_NET_0_74450, B => 
        HIEFFPLA_NET_0_74646, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74700);
    
    HIEFFPLA_INST_0_70702 : AND3
      port map(A => HIEFFPLA_NET_0_72034, B => 
        HIEFFPLA_NET_0_72033, C => \Timing_0/s_time[4]_net_1\, Y
         => HIEFFPLA_NET_0_72038);
    
    HIEFFPLA_INST_0_58083 : AO1
      port map(A => \Sensors_0_gyro_y[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75155, Y => HIEFFPLA_NET_0_74859);
    
    \General_Controller_0/status_bits_1[50]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74196, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[50]\);
    
    HIEFFPLA_INST_0_63098 : NAND3C
      port map(A => HIEFFPLA_NET_0_73828, B => 
        HIEFFPLA_NET_0_73850, C => HIEFFPLA_NET_0_74024, Y => 
        HIEFFPLA_NET_0_73829);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[8]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72553, Q => 
        \Sensors_0_gyro_x[8]\);
    
    HIEFFPLA_INST_0_64116 : OR2A
      port map(A => HIEFFPLA_NET_0_73579, B => 
        \General_Controller_0/constant_bias_voltage_0[15]_net_1\, 
        Y => HIEFFPLA_NET_0_73666);
    
    HIEFFPLA_INST_0_54932 : NOR2A
      port map(A => \ClockDivs_0/cnt_800kHz[1]_net_1\, B => 
        \ClockDivs_0/cnt_800kHz[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75636);
    
    HIEFFPLA_INST_0_66774 : AO1
      port map(A => HIEFFPLA_NET_0_73055, B => 
        HIEFFPLA_NET_0_73097, C => HIEFFPLA_NET_0_73028, Y => 
        HIEFFPLA_NET_0_73037);
    
    HIEFFPLA_INST_0_57159 : AND2
      port map(A => \Sensors_0_pressure_time[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, Y
         => HIEFFPLA_NET_0_75146);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_20\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[3]\\\\\, CLK => 
        CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_20_Q\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[0]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72482, Q => 
        \Sensors_0_gyro_y[0]\);
    
    HIEFFPLA_INST_0_69252 : NAND3C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, Y
         => HIEFFPLA_NET_0_72439);
    
    HIEFFPLA_INST_0_66115 : NAND2B
      port map(A => \Science_0/DAC_SET_0/state[2]_net_1\, B => 
        \Science_0/DAC_SET_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73205);
    
    HIEFFPLA_INST_0_55647 : NOR2A
      port map(A => HIEFFPLA_NET_0_75437, B => 
        \Communications_0/UART_1/rx_clk_count_c0\, Y => 
        HIEFFPLA_NET_0_75456);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[6]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75261, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\);
    
    HIEFFPLA_INST_0_70546 : NOR2A
      port map(A => \Timing_0/m_count[3]_net_1\, B => 
        \Timing_0/m_count[0]_net_1\, Y => HIEFFPLA_NET_0_72085);
    
    \Science_0/SET_LP_GAIN_0/old_G3[1]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73168, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/old_G3[1]_net_1\);
    
    HIEFFPLA_INST_0_69505 : MX2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[4]\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[6]\, 
        S => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72375);
    
    HIEFFPLA_INST_0_67344 : OR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72903);
    
    HIEFFPLA_INST_0_56499 : AX1
      port map(A => HIEFFPLA_NET_0_75350, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, C
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, 
        Y => HIEFFPLA_NET_0_75263);
    
    HIEFFPLA_INST_0_59431 : MX2A
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        HIEFFPLA_NET_0_74486, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74555);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[22]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[22]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[22]\);
    
    HIEFFPLA_INST_0_70032 : NAND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72241);
    
    HIEFFPLA_INST_0_66070 : AX1C
      port map(A => \Science_0/DAC_SET_0/cnt[0]_net_1\, B => 
        HIEFFPLA_NET_0_73213, C => 
        \Science_0/DAC_SET_0/cnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73218);
    
    HIEFFPLA_INST_0_57756 : AOI1
      port map(A => \Science_0_exp_packet_0[50]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74816, Y => HIEFFPLA_NET_0_74952);
    
    \General_Controller_0/en_science_packets\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74315, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74314, Q => 
        General_Controller_0_en_science_packets);
    
    \Data_Saving_0/Packet_Saver_0/data_out[19]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75226, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[19]\);
    
    HIEFFPLA_INST_0_63344 : MX2
      port map(A => HIEFFPLA_NET_0_74127, B => 
        HIEFFPLA_NET_0_73537, S => HIEFFPLA_NET_0_73965, Y => 
        HIEFFPLA_NET_0_73773);
    
    \General_Controller_0/constant_bias_voltage_0[8]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[8]_net_1\);
    
    \L3WR_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => L3WR_c, E => \VCC\, DOUT => 
        \L3WR_pad/U0/NET1\, EOUT => \L3WR_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_65702 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt4up[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt4up[0]_net_1\, C => 
        HIEFFPLA_NET_0_73309, Y => HIEFFPLA_NET_0_73305);
    
    HIEFFPLA_INST_0_57167 : AO1
      port map(A => \Sensors_0_gyro_time[18]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75141, Y => HIEFFPLA_NET_0_75142);
    
    \Science_0/ADC_READ_0/exp_packet_1[51]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[17]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[51]\);
    
    HIEFFPLA_INST_0_61127 : AO1A
      port map(A => HIEFFPLA_NET_0_74327, B => 
        HIEFFPLA_NET_0_74333, C => HIEFFPLA_NET_0_74269, Y => 
        HIEFFPLA_NET_0_74270);
    
    HIEFFPLA_INST_0_57285 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[45]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75095);
    
    AFLSDF_INV_35 : INV
      port map(A => HIEFFPLA_NET_0_72277, Y => \AFLSDF_INV_35\);
    
    \Science_0/ADC_READ_0/chan3_data[4]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[4]\);
    
    HIEFFPLA_INST_0_67077 : AOI1C
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        B => HIEFFPLA_NET_0_72739, C => HIEFFPLA_NET_0_72929, Y
         => HIEFFPLA_NET_0_72970);
    
    HIEFFPLA_INST_0_66647 : AND3
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_net_1\, B
         => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_1_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_2_net_1\, 
        Y => sda_cl_1_RNIBFPP);
    
    \General_Controller_0/sweep_table_samples_per_point[9]\ : 
        DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[9]_net_1\);
    
    \General_Controller_0/constant_bias_voltage_1[14]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[14]_net_1\);
    
    \General_Controller_0/constant_bias_voltage_1[12]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[12]_net_1\);
    
    HIEFFPLA_INST_0_69536 : AO1A
      port map(A => HIEFFPLA_NET_0_72364, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        C => \Sensors_0/Pressure_Sensor_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72369);
    
    \General_Controller_0/uc_tx_nextstate[6]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73623, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73857, Q => 
        \General_Controller_0/uc_tx_nextstate[6]_net_1\);
    
    \General_Controller_0/st_raddr[7]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[7]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73979, Q => 
        \General_Controller_0_st_raddr_1[7]\);
    
    HIEFFPLA_INST_0_57496 : AND2
      port map(A => \Science_0_exp_packet_0[19]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, Y
         => HIEFFPLA_NET_0_75029);
    
    \General_Controller_0/state_seconds[12]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74237, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[12]_net_1\);
    
    \Timing_0/m_count[5]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72074, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_count[5]_net_1\);
    
    HIEFFPLA_INST_0_62416 : AO1A
      port map(A => HIEFFPLA_NET_0_74080, B => 
        HIEFFPLA_NET_0_74085, C => HIEFFPLA_NET_0_74103, Y => 
        HIEFFPLA_NET_0_73986);
    
    \Timing_0/f_time[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72088, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/f_time[2]_net_1\);
    
    HIEFFPLA_INST_0_57724 : NAND3C
      port map(A => HIEFFPLA_NET_0_74843, B => 
        HIEFFPLA_NET_0_74834, C => HIEFFPLA_NET_0_74820, Y => 
        HIEFFPLA_NET_0_74959);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[6]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[6]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[6]\);
    
    \Communications_0/UART_0/tx_clk_count[8]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75518, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_clk_count_i_0[8]\);
    
    HIEFFPLA_INST_0_59197 : AND3B
      port map(A => HIEFFPLA_NET_0_74344, B => 
        Communications_0_ext_tx_rdy, C => 
        \GS_Readout_0/state[5]_net_1\, Y => HIEFFPLA_NET_0_74590);
    
    HIEFFPLA_INST_0_65358 : XA1B
      port map(A => HIEFFPLA_NET_0_73399, B => 
        \Science_0/ADC_READ_0/cnt1dn[7]_net_1\, C => 
        HIEFFPLA_NET_0_73244, Y => HIEFFPLA_NET_0_73401);
    
    HIEFFPLA_INST_0_61828 : NAND2B
      port map(A => UC_PWR_EN_c, B => 
        \General_Controller_0/flight_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74120);
    
    HIEFFPLA_INST_0_63279 : NOR2A
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_substate[0]_net_1\, Y
         => HIEFFPLA_NET_0_73791);
    
    HIEFFPLA_INST_0_57857 : AO1B
      port map(A => \Sensors_0_mag_time[21]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74923, Y => HIEFFPLA_NET_0_74924);
    
    \General_Controller_0/sweep_table_sample_skip[15]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[15]_net_1\);
    
    HIEFFPLA_INST_0_69122 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[3]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[4]_net_1\, 
        C => HIEFFPLA_NET_0_72557, Y => HIEFFPLA_NET_0_72466);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[3]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72276, Q => \Sensors_0_pressure_raw[3]\);
    
    HIEFFPLA_INST_0_65035 : XA1
      port map(A => HIEFFPLA_NET_0_73448, B => 
        \Pressure_Signal_Debounce_0/ms_cnt[9]_net_1\, C => 
        HIEFFPLA_NET_0_73477, Y => HIEFFPLA_NET_0_73484);
    
    HIEFFPLA_INST_0_65176 : AOI1
      port map(A => HIEFFPLA_NET_0_73463, B => 
        \Sensors_0_pressure_raw[22]\, C => 
        \Sensors_0_pressure_raw[23]\, Y => HIEFFPLA_NET_0_73452);
    
    HIEFFPLA_INST_0_61600 : AND3
      port map(A => HIEFFPLA_NET_0_73778, B => 
        HIEFFPLA_NET_0_74172, C => HIEFFPLA_NET_0_73972, Y => 
        HIEFFPLA_NET_0_74176);
    
    HIEFFPLA_INST_0_64589 : NOR3B
      port map(A => \General_Controller_0/uc_tx_state[7]_net_1\, 
        B => HIEFFPLA_NET_0_74319, C => HIEFFPLA_NET_0_74324, Y
         => HIEFFPLA_NET_0_73594);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/temp[4]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72555, Q => 
        \Sensors_0_gyro_temp[4]\);
    
    HIEFFPLA_INST_0_59857 : AND2
      port map(A => HIEFFPLA_NET_0_74448, B => 
        HIEFFPLA_NET_0_74397, Y => HIEFFPLA_NET_0_74496);
    
    \Science_0/ADC_READ_0/exp_packet_1[49]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[15]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[49]\);
    
    HIEFFPLA_INST_0_69138 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[7]_net_1\, 
        C => HIEFFPLA_NET_0_72557, Y => HIEFFPLA_NET_0_72462);
    
    HIEFFPLA_INST_0_57030 : MX2
      port map(A => HIEFFPLA_NET_0_75038, B => 
        HIEFFPLA_NET_0_74955, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75179);
    
    HIEFFPLA_INST_0_71011 : MX2C
      port map(A => HIEFFPLA_NET_0_73506, B => 
        HIEFFPLA_NET_0_73518, S => 
        \I2C_PassThrough_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_71990);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[1]\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_73129, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73041, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[1]_net_1\);
    
    HIEFFPLA_INST_0_60153 : MX2
      port map(A => \Science_0_chan5_data[1]\, B => 
        \Science_0_chan5_data[5]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74453);
    
    \General_Controller_0/sweep_table_probe_id[5]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73924, Q => 
        \General_Controller_0/sweep_table_probe_id[5]_net_1\);
    
    HIEFFPLA_INST_0_55026 : AND3
      port map(A => HIEFFPLA_NET_0_75593, B => 
        HIEFFPLA_NET_0_75591, C => HIEFFPLA_NET_0_75602, Y => 
        HIEFFPLA_NET_0_75611);
    
    HIEFFPLA_INST_0_55865 : NAND2B
      port map(A => HIEFFPLA_NET_0_75400, B => 
        HIEFFPLA_NET_0_75419, Y => HIEFFPLA_NET_0_75409);
    
    \I2C_PassThrough_0/state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73513, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \I2C_PassThrough_0/state[0]_net_1\);
    
    \Science_0/SET_LP_GAIN_0/old_G1[1]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73176, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/old_G1[1]_net_1\);
    
    \Communications_0/UART_1/rx_byte[1]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75378, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75495, Q => 
        \Communications_0/UART_1/rx_byte[1]_net_1\);
    
    HIEFFPLA_INST_0_66609 : MX2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[3]\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_data_out[7]\, 
        S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73084);
    
    HIEFFPLA_INST_0_64773 : NOR3B
      port map(A => HIEFFPLA_NET_0_73592, B => 
        HIEFFPLA_NET_0_73543, C => 
        \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73544);
    
    HIEFFPLA_INST_0_62320 : NAND2B
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74006);
    
    \Science_0/ADC_READ_0/cnt3up[2]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73334, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3up[2]_net_1\);
    
    HIEFFPLA_INST_0_59707 : AO1
      port map(A => HIEFFPLA_NET_0_74420, B => 
        HIEFFPLA_NET_0_74341, C => HIEFFPLA_NET_0_74400, Y => 
        HIEFFPLA_NET_0_74519);
    
    HIEFFPLA_INST_0_65063 : OA1C
      port map(A => HIEFFPLA_NET_0_73479, B => 
        \Pressure_Signal_Debounce_0/state[0]_net_1\, C => 
        CLKINT_1_Y, Y => HIEFFPLA_NET_0_73478);
    
    HIEFFPLA_INST_0_56551 : NOR2A
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[9]_net_1\, B
         => \Data_Saving_0/FPGA_Buffer_0_afull\, Y => 
        HIEFFPLA_NET_0_75242);
    
    HIEFFPLA_INST_0_64557 : AO1A
      port map(A => HIEFFPLA_NET_0_73556, B => 
        HIEFFPLA_NET_0_73577, C => HIEFFPLA_NET_0_73581, Y => 
        HIEFFPLA_NET_0_73601);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[10]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72807, Q => 
        \Sensors_0_mag_z[10]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[10]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72777, Q => 
        \Sensors_0_acc_y[10]\);
    
    HIEFFPLA_INST_0_60011 : NOR2A
      port map(A => HIEFFPLA_NET_0_74410, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74474);
    
    HIEFFPLA_INST_0_70518 : XOR2
      port map(A => HIEFFPLA_NET_0_72125, B => 
        \Timekeeper_0_milliseconds[3]\, Y => HIEFFPLA_NET_0_72099);
    
    HIEFFPLA_INST_0_61577 : OR3A
      port map(A => HIEFFPLA_NET_0_74182, B => 
        \General_Controller_0/sweep_table_probe_id[4]_net_1\, C
         => \General_Controller_0/sweep_table_probe_id[5]_net_1\, 
        Y => HIEFFPLA_NET_0_74180);
    
    HIEFFPLA_INST_0_55615 : XA1
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\, B => 
        HIEFFPLA_NET_0_75477, C => HIEFFPLA_NET_0_75437, Y => 
        HIEFFPLA_NET_0_75464);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[5]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72489, Q => 
        \ch3_data_net_0[1]\);
    
    HIEFFPLA_INST_0_69264 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, C
         => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72434);
    
    \FMC_DA_pad[7]/U0/U0\ : IOPAD_TRI
      port map(D => \FMC_DA_pad[7]/U0/NET1\, E => 
        \FMC_DA_pad[7]/U0/NET2\, PAD => FMC_DA(7));
    
    \General_Controller_0/constant_bias_voltage_1[0]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[0]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[0]_net_1\);
    
    \TOP_UART_RX_pad/U0/U1\ : IOIN_IB
      port map(YIN => \TOP_UART_RX_pad/U0/NET1\, Y => 
        TOP_UART_RX_c);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[3]\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_73127, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73041, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[3]_net_1\);
    
    HIEFFPLA_INST_0_65439 : XA1B
      port map(A => \Science_0/ADC_READ_0/cnt2dn[0]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2dn[1]_net_1\, C => 
        HIEFFPLA_NET_0_73381, Y => HIEFFPLA_NET_0_73375);
    
    HIEFFPLA_INST_0_68611 : AOI1
      port map(A => \Sensors_0/Gyro_0/L3GD20H_Interface_0_we\, B
         => \Sensors_0/Gyro_0/state[8]\, C => 
        HIEFFPLA_NET_0_72605, Y => HIEFFPLA_NET_0_72606);
    
    HIEFFPLA_INST_0_68447 : AO1
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[2]_net_1\, B => 
        GYRO_SCL_c, C => HIEFFPLA_NET_0_72621, Y => 
        HIEFFPLA_NET_0_72648);
    
    \General_Controller_0/temp_first_byte[4]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73872, Q => 
        \General_Controller_0/temp_first_byte[4]_net_1\);
    
    HIEFFPLA_INST_0_65630 : AND2
      port map(A => \Science_0/ADC_READ_0/cnt4dn[0]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt4dn[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73324);
    
    HIEFFPLA_INST_0_69470 : NOR3B
      port map(A => HIEFFPLA_NET_0_72410, B => 
        HIEFFPLA_NET_0_72346, C => PRESSURE_SCL_c, Y => 
        HIEFFPLA_NET_0_72381);
    
    HIEFFPLA_INST_0_69313 : AO1A
      port map(A => HIEFFPLA_NET_0_72344, B => 
        HIEFFPLA_NET_0_72419, C => HIEFFPLA_NET_0_72420, Y => 
        HIEFFPLA_NET_0_72421);
    
    HIEFFPLA_INST_0_66922 : AO1
      port map(A => HIEFFPLA_NET_0_72762, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        C => HIEFFPLA_NET_0_72751, Y => HIEFFPLA_NET_0_73004);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_7\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[7]\\\\\, CLK => 
        CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_7_Q\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73032, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\);
    
    HIEFFPLA_INST_0_61711 : MX2
      port map(A => \SweepTable_0_RD[8]\, B => 
        \SweepTable_1_RD[8]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74156);
    
    HIEFFPLA_INST_0_57982 : AO1
      port map(A => \Science_0_exp_packet_0[30]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74785, Y => HIEFFPLA_NET_0_74888);
    
    \Communications_0/UART_1/rx_byte[3]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75378, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75493, Q => 
        \Communications_0/UART_1/rx_byte[3]_net_1\);
    
    HIEFFPLA_INST_0_65281 : OR3A
      port map(A => \Science_0/ADC_READ_0/chan[0]_net_1\, B => 
        \Science_0/ADC_READ_0/chan[1]_net_1\, C => 
        HIEFFPLA_NET_0_73243, Y => HIEFFPLA_NET_0_73424);
    
    HIEFFPLA_INST_0_59019 : NAND3B
      port map(A => \GS_Readout_0/state[1]_net_1\, B => 
        \GS_Readout_0/state[2]_net_1\, C => HIEFFPLA_NET_0_74635, 
        Y => HIEFFPLA_NET_0_74636);
    
    HIEFFPLA_INST_0_57136 : AND2
      port map(A => \Sensors_0_pressure_temp_raw[16]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75161);
    
    HIEFFPLA_INST_0_61380 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[40]\, B => 
        \Timekeeper_0_milliseconds[0]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74206);
    
    HIEFFPLA_INST_0_57231 : AO1
      port map(A => \Sensors_0_pressure_time[17]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75080, Y => HIEFFPLA_NET_0_75119);
    
    HIEFFPLA_INST_0_56682 : MX2
      port map(A => HIEFFPLA_NET_0_75192, B => 
        HIEFFPLA_NET_0_75054, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75225);
    
    HIEFFPLA_INST_0_62252 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state_0[1]_net_1\, 
        B => \General_Controller_0/uc_rx_substate[2]_net_1\, C
         => HIEFFPLA_NET_0_73810, Y => HIEFFPLA_NET_0_74020);
    
    HIEFFPLA_INST_0_70401 : XOR2
      port map(A => HIEFFPLA_NET_0_72155, B => 
        \Timekeeper_0_microseconds[13]\, Y => 
        HIEFFPLA_NET_0_72147);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRY[8]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75295, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[8]\\\\\);
    
    \Timekeeper_0/milliseconds[18]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72107, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[18]\);
    
    \GS_Readout_0/prevState[4]\ : DFN1E0C1
      port map(D => \GS_Readout_0/state[4]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \GS_Readout_0/state[6]_net_1\, Q => 
        \GS_Readout_0/prevState[4]_net_1\);
    
    HIEFFPLA_INST_0_60659 : MX2
      port map(A => HIEFFPLA_NET_0_74401, B => 
        HIEFFPLA_NET_0_74513, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74380);
    
    HIEFFPLA_INST_0_55988 : AND2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\, B
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, 
        Y => HIEFFPLA_NET_0_75376);
    
    HIEFFPLA_INST_0_70513 : AX1C
      port map(A => \Timekeeper_0_milliseconds[22]\, B => 
        HIEFFPLA_NET_0_72122, C => 
        \Timekeeper_0_milliseconds[23]\, Y => 
        HIEFFPLA_NET_0_72101);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[7]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72462, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[7]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[15]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72490, Q => 
        \ch3_data_net_0[11]\);
    
    HIEFFPLA_INST_0_56546 : AX1
      port map(A => HIEFFPLA_NET_0_75243, B => 
        \Data_Saving_0/Interrupt_Generator_0/counter[7]_net_1\, C
         => 
        \Data_Saving_0/Interrupt_Generator_0/counter[9]_net_1\, Y
         => HIEFFPLA_NET_0_75244);
    
    HIEFFPLA_INST_0_64821 : AND3B
      port map(A => HIEFFPLA_NET_0_73523, B => 
        HIEFFPLA_NET_0_73526, C => 
        \General_Controller_0/uc_tx_substate[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73532);
    
    HIEFFPLA_INST_0_59863 : MX2
      port map(A => \Sensors_0_pressure_temp_raw[23]\, B => 
        \Sensors_0_pressure_raw[15]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74495);
    
    HIEFFPLA_INST_0_56542 : AX1C
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[7]_net_1\, B
         => HIEFFPLA_NET_0_75255, C => 
        \Data_Saving_0/Interrupt_Generator_0/counter[8]_net_1\, Y
         => HIEFFPLA_NET_0_75245);
    
    \Science_0/DAC_SET_0/vector[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73186, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[0]_net_1\);
    
    HIEFFPLA_INST_0_62574 : NAND3C
      port map(A => HIEFFPLA_NET_0_73980, B => 
        HIEFFPLA_NET_0_73967, C => HIEFFPLA_NET_0_73932, Y => 
        HIEFFPLA_NET_0_73953);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[6]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72777, Q => 
        \Sensors_0_acc_y[6]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[3]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72865, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[3]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[28]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[12]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[28]\);
    
    HIEFFPLA_INST_0_56148 : AO13
      port map(A => HIEFFPLA_NET_0_75294, B => 
        HIEFFPLA_NET_0_75275, C => HIEFFPLA_NET_0_75279, Y => 
        HIEFFPLA_NET_0_75339);
    
    HIEFFPLA_INST_0_68054 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72743);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[4]\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72296, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72221, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[4]_net_1\);
    
    \Science_0/DAC_SET_0/vector[12]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73201, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[12]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[4]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72808, Q => 
        \Sensors_0_mag_z[4]\);
    
    HIEFFPLA_INST_0_59615 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[2]\, B => 
        \Data_Hub_Packets_0_status_packet[6]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74531);
    
    HIEFFPLA_INST_0_57154 : AND2
      port map(A => \Sensors_0_pressure_time[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, Y
         => HIEFFPLA_NET_0_75151);
    
    \Science_0/ADC_READ_0/chan1_data[5]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[5]\);
    
    \General_Controller_0/constant_bias_voltage_0[15]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[15]_net_1\);
    
    \Science_0/ADC_READ_0/cnt4up[0]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73306, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4up[0]_net_1\);
    
    HIEFFPLA_INST_0_64327 : MX2
      port map(A => HIEFFPLA_NET_0_73725, B => 
        HIEFFPLA_NET_0_73717, S => HIEFFPLA_NET_0_73619, Y => 
        HIEFFPLA_NET_0_73637);
    
    HIEFFPLA_INST_0_59154 : AND3C
      port map(A => HIEFFPLA_NET_0_74595, B => 
        HIEFFPLA_NET_0_74589, C => HIEFFPLA_NET_0_74583, Y => 
        HIEFFPLA_NET_0_74599);
    
    HIEFFPLA_INST_0_68000 : NAND2B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72756);
    
    \Communications_0/UART_0/rx_clk_count[28]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75571, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75554, Q => 
        \Communications_0/UART_0/rx_clk_count[28]_net_1\);
    
    HIEFFPLA_INST_0_63092 : NAND3
      port map(A => HIEFFPLA_NET_0_74091, B => 
        HIEFFPLA_NET_0_73842, C => HIEFFPLA_NET_0_73803, Y => 
        HIEFFPLA_NET_0_73830);
    
    HIEFFPLA_INST_0_61895 : AND2
      port map(A => \General_Controller_0/uc_rx_byte[2]_net_1\, B
         => \General_Controller_0/uc_rx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74105);
    
    HIEFFPLA_INST_0_67218 : AND3
      port map(A => HIEFFPLA_NET_0_72949, B => 
        HIEFFPLA_NET_0_72950, C => HIEFFPLA_NET_0_72957, Y => 
        HIEFFPLA_NET_0_72936);
    
    HIEFFPLA_INST_0_63842 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[3]_net_1\, B
         => 
        \General_Controller_0/sweep_table_sample_skip[3]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73702);
    
    HIEFFPLA_INST_0_70377 : AND3
      port map(A => \Timekeeper_0_microseconds[3]\, B => 
        HIEFFPLA_NET_0_72154, C => \Timekeeper_0_microseconds[4]\, 
        Y => HIEFFPLA_NET_0_72156);
    
    \Science_0/ADC_READ_0/cnt3dn[0]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73347, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3dn[0]_net_1\);
    
    HIEFFPLA_INST_0_58591 : NOR3B
      port map(A => \Eject_Signal_Debounce_0/ms_cnt[4]_net_1\, B
         => \Eject_Signal_Debounce_0/ms_cnt[2]_net_1\, C => 
        HIEFFPLA_NET_0_74726, Y => HIEFFPLA_NET_0_74727);
    
    HIEFFPLA_INST_0_57870 : AOI1
      port map(A => \Sensors_0_acc_time[22]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74919, Y => HIEFFPLA_NET_0_74920);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[9]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72490, Q => 
        \ch3_data_net_0[5]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[11]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[11]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[11]\);
    
    HIEFFPLA_INST_0_69754 : OA1C
      port map(A => \Sensors_0/Pressure_Sensor_0/state[8]\, B => 
        HIEFFPLA_NET_0_72285, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72315);
    
    HIEFFPLA_INST_0_64157 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_1[5]_net_1\, 
        B => 
        \General_Controller_0/constant_bias_voltage_1[13]_net_1\, 
        S => \General_Controller_0/uc_tx_substate[1]_net_1\, Y
         => HIEFFPLA_NET_0_73660);
    
    \Science_0/ADC_READ_0/exp_packet_1[66]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[10]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[66]\);
    
    HIEFFPLA_INST_0_68174 : NOR3B
      port map(A => HIEFFPLA_NET_0_72772, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        C => HIEFFPLA_NET_0_72902, Y => HIEFFPLA_NET_0_72716);
    
    \General_Controller_0/constant_bias_probe_id[1]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73923, Q => 
        \General_Controller_0/un10_uc_tx_rdy_i[1]\);
    
    HIEFFPLA_INST_0_68383 : AND2B
      port map(A => \Sensors_0/Gyro_0/state[8]\, B => GYRO_SCL_c, 
        Y => HIEFFPLA_NET_0_72662);
    
    HIEFFPLA_INST_0_67057 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[2]\, 
        B => \Sensors_0/Accelerometer_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72976);
    
    \General_Controller_0/sweep_table_sweep_cnt[14]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74139, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[14]_net_1\);
    
    \Science_0/DAC_SET_0/vector[13]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73200, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[13]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[20]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[4]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[20]\);
    
    HIEFFPLA_INST_0_66021 : AX1C
      port map(A => \Science_0/ADC_READ_0/cnt_chan[0]_net_1\, B
         => HIEFFPLA_NET_0_73241, C => 
        \Science_0/ADC_READ_0/cnt_chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73236);
    
    HIEFFPLA_INST_0_60561 : MX2
      port map(A => HIEFFPLA_NET_0_74542, B => 
        HIEFFPLA_NET_0_74389, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74395);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[7]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[7]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[7]\);
    
    HIEFFPLA_INST_0_57004 : MX2
      port map(A => HIEFFPLA_NET_0_75045, B => 
        HIEFFPLA_NET_0_74959, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75183);
    
    HIEFFPLA_INST_0_58361 : AO1
      port map(A => \Sensors_0_acc_y[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74791, Y => HIEFFPLA_NET_0_74792);
    
    HIEFFPLA_INST_0_57995 : AO1
      port map(A => \Science_0_exp_packet_0[54]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_74811, Y => HIEFFPLA_NET_0_74884);
    
    \Timekeeper_0/microseconds[14]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72146, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[14]\);
    
    \General_Controller_0/constant_bias_voltage_0[0]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[0]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[0]_net_1\);
    
    \Timing_0/m_count[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72077, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_count[3]_net_1\);
    
    \ClockDivs_0/cnt_800kHz[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75634, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \ClockDivs_0/cnt_800kHz[2]_net_1\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/state_0[8]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73061, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/state_0[8]\);
    
    HIEFFPLA_INST_0_64020 : MX2
      port map(A => HIEFFPLA_NET_0_73650, B => 
        HIEFFPLA_NET_0_73642, S => HIEFFPLA_NET_0_73599, Y => 
        HIEFFPLA_NET_0_73679);
    
    HIEFFPLA_INST_0_59743 : MX2
      port map(A => HIEFFPLA_NET_0_74413, B => 
        HIEFFPLA_NET_0_74406, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74514);
    
    HIEFFPLA_INST_0_69050 : AND3
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        B => \Sensors_0/Gyro_0/state[8]\, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, Y
         => HIEFFPLA_NET_0_72485);
    
    \Communications_0/FFU_Command_Checker_0/command_out[4]\ : 
        DFN1E1C1
      port map(D => \Communications_0/UART_0_recv[4]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75625, Q => \Communications_0_ext_recv[4]\);
    
    HIEFFPLA_INST_0_70079 : OR3B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[3]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72227);
    
    \Data_Saving_0/Packet_Saver_0/data_out[21]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75223, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[21]\);
    
    HIEFFPLA_INST_0_60814 : XA1B
      port map(A => \GS_Readout_0/subState[1]_net_1\, B => 
        HIEFFPLA_NET_0_74348, C => HIEFFPLA_NET_0_74350, Y => 
        HIEFFPLA_NET_0_74354);
    
    HIEFFPLA_INST_0_62391 : AOI5
      port map(A => HIEFFPLA_NET_0_73811, B => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73991);
    
    HIEFFPLA_INST_0_63554 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[11]_net_1\, B
         => \General_Controller_0/sweep_table_points[11]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73750);
    
    HIEFFPLA_INST_0_56063 : XA1A
      port map(A => HIEFFPLA_NET_0_75263, B => 
        HIEFFPLA_NET_0_75270, C => HIEFFPLA_NET_0_75325, Y => 
        HIEFFPLA_NET_0_75357);
    
    \General_Controller_0/status_bits_1[54]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74192, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[54]\);
    
    HIEFFPLA_INST_0_68365 : AND2
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, B
         => HIEFFPLA_NET_0_72689, Y => HIEFFPLA_NET_0_72670);
    
    HIEFFPLA_INST_0_65719 : AND2
      port map(A => \Science_0/ADC_READ_0/cnt4up[3]_net_1\, B => 
        HIEFFPLA_NET_0_73307, Y => HIEFFPLA_NET_0_73300);
    
    HIEFFPLA_INST_0_64602 : AND3C
      port map(A => \General_Controller_0/uc_tx_state[5]_net_1\, 
        B => \General_Controller_0/uc_tx_state[1]_net_1\, C => 
        \General_Controller_0/uc_tx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73591);
    
    HIEFFPLA_INST_0_59763 : MX2
      port map(A => \Sensors_0_pressure_temp_raw[22]\, B => 
        \Sensors_0_pressure_raw[14]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74512);
    
    \General_Controller_0/uc_tx_substate[4]\ : DFN1C1
      port map(D => 
        \General_Controller_0/uc_tx_substate[4]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_tx_substate[4]_net_1\);
    
    HIEFFPLA_INST_0_64525 : AO1A
      port map(A => HIEFFPLA_NET_0_73556, B => 
        HIEFFPLA_NET_0_73615, C => HIEFFPLA_NET_0_73579, Y => 
        HIEFFPLA_NET_0_73607);
    
    HIEFFPLA_INST_0_63290 : OR3A
      port map(A => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[4]_net_1\, C => 
        \General_Controller_0/uc_rx_substate[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73786);
    
    HIEFFPLA_INST_0_61492 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[54]\, B => 
        \Timekeeper_0_milliseconds[14]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74192);
    
    HIEFFPLA_INST_0_70590 : AX1C
      port map(A => HIEFFPLA_NET_0_72068, B => 
        \Timing_0/m_time[6]_net_1\, C => \m_time[7]\, Y => 
        HIEFFPLA_NET_0_72071);
    
    HIEFFPLA_INST_0_58133 : AO1
      port map(A => \Sensors_0_mag_time[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75150, Y => HIEFFPLA_NET_0_74843);
    
    HIEFFPLA_INST_0_63782 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[1]_net_1\, 
        B => \General_Controller_0/sweep_table_points[1]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73712);
    
    HIEFFPLA_INST_0_68192 : AO1
      port map(A => HIEFFPLA_NET_0_72739, B => 
        \Sensors_0/Accelerometer_0/state_0[8]\, C => 
        HIEFFPLA_NET_0_72709, Y => HIEFFPLA_NET_0_72710);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[4]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72753, Q => 
        \Sensors_0_acc_z[4]\);
    
    HIEFFPLA_INST_0_70357 : AND3
      port map(A => \Timekeeper_0_microseconds[13]\, B => 
        HIEFFPLA_NET_0_72155, C => 
        \Timekeeper_0_microseconds[14]\, Y => 
        HIEFFPLA_NET_0_72161);
    
    \Communications_0/UART_0/rx_byte[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75380, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75605, Q => 
        \Communications_0/UART_0/rx_byte[7]_net_1\);
    
    HIEFFPLA_INST_0_71054 : AXO6
      port map(A => \General_Controller_0/uc_rx_byte[2]_net_1\, B
         => \General_Controller_0/uc_rx_byte[0]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[1]_net_1\, Y => 
        HIEFFPLA_NET_0_71985);
    
    HIEFFPLA_INST_0_69094 : NOR3A
      port map(A => HIEFFPLA_NET_0_72544, B => 
        HIEFFPLA_NET_0_72459, C => HIEFFPLA_NET_0_72453, Y => 
        HIEFFPLA_NET_0_72471);
    
    \Science_0/DAC_SET_0/ADR[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73229, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/ADR[0]_net_1\);
    
    HIEFFPLA_INST_0_58551 : XO1
      port map(A => FFU_EJECTED_c, B => 
        \Eject_Signal_Debounce_0/state[1]_net_1\, C => 
        \Eject_Signal_Debounce_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74737);
    
    HIEFFPLA_INST_0_65110 : AND3C
      port map(A => \Sensors_0_pressure_raw[2]\, B => 
        \Sensors_0_pressure_raw[0]\, C => 
        \Sensors_0_pressure_raw[3]\, Y => HIEFFPLA_NET_0_73469);
    
    \General_Controller_0/sweep_table_write_value[4]\ : DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[4]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[4]_net_1\);
    
    \General_Controller_0/sweep_table_samples_per_step[0]\ : 
        DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[0]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[0]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[11]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72753, Q => 
        \Sensors_0_acc_z[11]\);
    
    HIEFFPLA_INST_0_58492 : NAND3
      port map(A => \Eject_Signal_Debounce_0/ms_cnt[4]_net_1\, B
         => \Eject_Signal_Debounce_0/ms_cnt[5]_net_1\, C => 
        \Eject_Signal_Debounce_0/state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74750);
    
    HIEFFPLA_INST_0_68364 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, B => 
        HIEFFPLA_NET_0_72670, C => GYRO_SCL_c, Y => 
        HIEFFPLA_NET_0_72671);
    
    HIEFFPLA_INST_0_68148 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        Y => HIEFFPLA_NET_0_72722);
    
    HIEFFPLA_INST_0_61245 : XA1B
      port map(A => 
        \General_Controller_0/state_seconds[11]_net_1\, B => 
        HIEFFPLA_NET_0_74216, C => HIEFFPLA_NET_0_74217, Y => 
        HIEFFPLA_NET_0_74238);
    
    HIEFFPLA_INST_0_61182 : OA1C
      port map(A => \General_Controller_0/state_seconds[8]_net_1\, 
        B => HIEFFPLA_NET_0_74260, C => HIEFFPLA_NET_0_74259, Y
         => HIEFFPLA_NET_0_74257);
    
    HIEFFPLA_INST_0_59923 : MX2
      port map(A => HIEFFPLA_NET_0_74384, B => 
        HIEFFPLA_NET_0_74414, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74487);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/i2c_repeat_start\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72916, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72972, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_repeat_start\);
    
    HIEFFPLA_INST_0_62957 : AO1A
      port map(A => HIEFFPLA_NET_0_73886, B => 
        HIEFFPLA_NET_0_74103, C => HIEFFPLA_NET_0_73925, Y => 
        HIEFFPLA_NET_0_73858);
    
    HIEFFPLA_INST_0_58433 : NAND2B
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, B
         => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        Y => HIEFFPLA_NET_0_74768);
    
    HIEFFPLA_INST_0_59721 : NOR2A
      port map(A => HIEFFPLA_NET_0_74448, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74517);
    
    HIEFFPLA_INST_0_70059 : AO1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        B => HIEFFPLA_NET_0_72285, C => HIEFFPLA_NET_0_72224, Y
         => HIEFFPLA_NET_0_72232);
    
    HIEFFPLA_INST_0_69107 : OR3A
      port map(A => HIEFFPLA_NET_0_72544, B => 
        HIEFFPLA_NET_0_72457, C => HIEFFPLA_NET_0_72451, Y => 
        HIEFFPLA_NET_0_72469);
    
    \GS_Readout_0/state[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74609, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/state[2]_net_1\);
    
    \General_Controller_0/sweep_table_nof_steps[1]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73980, Q => 
        \General_Controller_0/sweep_table_nof_steps[1]_net_1\);
    
    HIEFFPLA_INST_0_55163 : XA1C
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[28]_net_1\, B => 
        HIEFFPLA_NET_0_75579, C => HIEFFPLA_NET_0_75567, Y => 
        HIEFFPLA_NET_0_75571);
    
    HIEFFPLA_INST_0_66026 : AND2B
      port map(A => \Science_0/ADC_RESET_0/state[0]_net_1\, B => 
        \Science_0/ADC_RESET_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73234);
    
    HIEFFPLA_INST_0_65239 : NOR3B
      port map(A => HIEFFPLA_NET_0_73433, B => 
        HIEFFPLA_NET_0_73436, C => \Sensors_0_pressure_raw[16]\, 
        Y => HIEFFPLA_NET_0_73437);
    
    HIEFFPLA_INST_0_68413 : MX2
      port map(A => HIEFFPLA_NET_0_72653, B => 
        HIEFFPLA_NET_0_72652, S => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_72656);
    
    HIEFFPLA_INST_0_57785 : AO1B
      port map(A => \Sensors_0_acc_x[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74942, Y => HIEFFPLA_NET_0_74943);
    
    HIEFFPLA_INST_0_67574 : AOI1C
      port map(A => HIEFFPLA_NET_0_72815, B => 
        HIEFFPLA_NET_0_72942, C => HIEFFPLA_NET_0_72914, Y => 
        HIEFFPLA_NET_0_72849);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[10]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72281, Q => \Sensors_0_pressure_raw[10]\);
    
    HIEFFPLA_INST_0_58699 : AO1
      port map(A => \General_Controller_0_gs_id[4]\, B => 
        HIEFFPLA_NET_0_74484, C => HIEFFPLA_NET_0_74645, Y => 
        HIEFFPLA_NET_0_74701);
    
    HIEFFPLA_INST_0_57923 : AO1
      port map(A => \Science_0_exp_packet_0[67]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75131, Y => HIEFFPLA_NET_0_74904);
    
    \Science_0/ADC_READ_0/chan2_data[6]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[6]\);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1P0_empty\ : DFN1P0
      port map(D => HIEFFPLA_NET_0_75368, CLK => CLKINT_2_Y, PRE
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/empty\);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_15\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[6]\\\\\, CLK => 
        CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_15_Q\);
    
    \Science_0/DAC_SET_0/state[4]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_73209, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/state[4]_net_1\);
    
    HIEFFPLA_INST_0_67448 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72877);
    
    \Communications_0/UART_0/tx_state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75499, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_state[1]_net_1\);
    
    HIEFFPLA_INST_0_65194 : AND3
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[8]_net_1\, 
        B => HIEFFPLA_NET_0_73444, C => HIEFFPLA_NET_0_73442, Y
         => HIEFFPLA_NET_0_73448);
    
    HIEFFPLA_INST_0_58354 : AO1
      port map(A => \Sensors_0_mag_y[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75105, Y => HIEFFPLA_NET_0_74794);
    
    HIEFFPLA_INST_0_65171 : AO1
      port map(A => HIEFFPLA_NET_0_73468, B => 
        HIEFFPLA_NET_0_73459, C => HIEFFPLA_NET_0_73452, Y => 
        HIEFFPLA_NET_0_73453);
    
    HIEFFPLA_INST_0_65210 : AND3
      port map(A => HIEFFPLA_NET_0_73444, B => 
        \Pressure_Signal_Debounce_0/ms_cnt[4]_net_1\, C => 
        \Pressure_Signal_Debounce_0/ms_cnt[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73445);
    
    AFLSDF_INV_31 : INV
      port map(A => CLKINT_1_Y, Y => \AFLSDF_INV_31\);
    
    \General_Controller_0/st_wdata[5]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[5]\);
    
    \Science_0/ADC_READ_0/state_0[1]\ : DFN1C1
      port map(D => \Science_0/ADC_READ_0/state[2]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, Q => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\);
    
    HIEFFPLA_INST_0_66536 : OR2A
      port map(A => HIEFFPLA_NET_0_73132, B => ACCE_SCL_c, Y => 
        HIEFFPLA_NET_0_73098);
    
    HIEFFPLA_INST_0_55500 : NOR3B
      port map(A => HIEFFPLA_NET_0_75487, B => 
        HIEFFPLA_NET_0_75488, C => 
        \Communications_0/UART_1/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75496);
    
    HIEFFPLA_INST_0_69284 : NOR3A
      port map(A => HIEFFPLA_NET_0_72348, B => 
        HIEFFPLA_NET_0_72426, C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72430);
    
    \Science_0/ADC_READ_0/exp_packet_1[4]\ : DFN1E0
      port map(D => \AFLSDF_INV_32\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[4]\);
    
    HIEFFPLA_INST_0_57795 : AO1B
      port map(A => \Sensors_0_gyro_x[13]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74939, Y => HIEFFPLA_NET_0_74940);
    
    HIEFFPLA_INST_0_55944 : XA1B
      port map(A => \Communications_0/UART_1/tx_state[1]_net_1\, 
        B => \Communications_0/UART_1/tx_state[0]_net_1\, C => 
        HIEFFPLA_NET_0_75420, Y => HIEFFPLA_NET_0_75388);
    
    \Communications_0/UART_0/rx_clk_count[23]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75576, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75554, Q => 
        \Communications_0/UART_0/rx_clk_count[23]_net_1\);
    
    HIEFFPLA_INST_0_57561 : AO1
      port map(A => \Sensors_0_pressure_raw[16]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_75007, Y => HIEFFPLA_NET_0_75008);
    
    HIEFFPLA_INST_0_55769 : AXO5
      port map(A => HIEFFPLA_NET_0_75427, B => 
        \Communications_0/UART_1/tx_state[1]_net_1\, C => 
        \Communications_0/UART_1/tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75428);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_14\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[3]\\\\\, CLK => 
        CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_14_Q\);
    
    HIEFFPLA_INST_0_55906 : AX1B
      port map(A => HIEFFPLA_NET_0_75386, B => 
        HIEFFPLA_NET_0_75417, C => 
        \Communications_0/UART_1/tx_clk_count_i_0[2]\, Y => 
        HIEFFPLA_NET_0_75400);
    
    HIEFFPLA_INST_0_69783 : AND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72306);
    
    HIEFFPLA_INST_0_68780 : AO1B
      port map(A => HIEFFPLA_NET_0_72563, B => 
        Sensors_0_gyro_new_data, C => HIEFFPLA_NET_0_72479, Y => 
        HIEFFPLA_NET_0_72564);
    
    HIEFFPLA_INST_0_65540 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt3dn[2]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt3dn[1]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt3dn[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73348);
    
    HIEFFPLA_INST_0_65895 : NAND3
      port map(A => \Science_0/ADC_READ_0_G1[0]\, B => 
        \Science_0/ADC_READ_0/cnt1up[4]_net_1\, C => 
        HIEFFPLA_NET_0_73276, Y => HIEFFPLA_NET_0_73262);
    
    HIEFFPLA_INST_0_60998 : NOR3A
      port map(A => HIEFFPLA_NET_0_74301, B => 
        \General_Controller_0/ext_rx_state[0]_net_1\, C => 
        CLKINT_1_Y, Y => HIEFFPLA_NET_0_74300);
    
    \General_Controller_0/status_bits_1[48]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74198, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[48]\);
    
    HIEFFPLA_INST_0_65448 : XA1C
      port map(A => \Science_0/ADC_READ_0/cnt2dn[3]_net_1\, B => 
        HIEFFPLA_NET_0_73377, C => HIEFFPLA_NET_0_73381, Y => 
        HIEFFPLA_NET_0_73373);
    
    HIEFFPLA_INST_0_62328 : AND3C
      port map(A => HIEFFPLA_NET_0_74003, B => 
        HIEFFPLA_NET_0_73909, C => 
        \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74004);
    
    HIEFFPLA_INST_0_70743 : AND3
      port map(A => \Timing_0/s_count[2]_net_1\, B => 
        HIEFFPLA_NET_0_72026, C => \Timing_0/s_count[1]_net_1\, Y
         => HIEFFPLA_NET_0_72025);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[5]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72919, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[5]_net_1\);
    
    \General_Controller_0/uc_rx_state_0[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74065, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\);
    
    HIEFFPLA_INST_0_57850 : AOI1
      port map(A => \Sensors_0_acc_time[20]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74925, Y => HIEFFPLA_NET_0_74926);
    
    HIEFFPLA_INST_0_65772 : AX1C
      port map(A => \Science_0/ADC_READ_0/cnt[5]_net_1\, B => 
        HIEFFPLA_NET_0_73293, C => 
        \Science_0/ADC_READ_0/cnt[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73283);
    
    HIEFFPLA_INST_0_65665 : XA1
      port map(A => HIEFFPLA_NET_0_73326, B => 
        \Science_0/ADC_READ_0/cnt4dn[4]_net_1\, C => 
        HIEFFPLA_NET_0_73274, Y => HIEFFPLA_NET_0_73314);
    
    HIEFFPLA_INST_0_65631 : AND2B
      port map(A => \Science_0/ADC_READ_0/cnt4dn[2]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt4dn[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73323);
    
    HIEFFPLA_INST_0_64995 : XA1
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[2]_net_1\, 
        B => HIEFFPLA_NET_0_73443, C => HIEFFPLA_NET_0_73490, Y
         => HIEFFPLA_NET_0_73493);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/temp[3]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72555, Q => 
        \Sensors_0_gyro_temp[3]\);
    
    \General_Controller_0/sweep_table_write_value[1]\ : DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[1]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[1]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_WADDR[2]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75312, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[2]\\\\\);
    
    HIEFFPLA_INST_0_62581 : OA1A
      port map(A => HIEFFPLA_NET_0_73897, B => 
        HIEFFPLA_NET_0_74037, C => HIEFFPLA_NET_0_73937, Y => 
        HIEFFPLA_NET_0_73952);
    
    HIEFFPLA_INST_0_61266 : AND2A
      port map(A => HIEFFPLA_NET_0_74217, B => 
        HIEFFPLA_NET_0_74231, Y => HIEFFPLA_NET_0_74232);
    
    HIEFFPLA_INST_0_57806 : AO1
      port map(A => \Sensors_0_mag_x[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74779, Y => HIEFFPLA_NET_0_74937);
    
    \Science_0/ADC_READ_0/exp_packet_1[64]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[8]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[64]\);
    
    HIEFFPLA_INST_0_62235 : AND3
      port map(A => HIEFFPLA_NET_0_73896, B => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, C => 
        HIEFFPLA_NET_0_73780, Y => HIEFFPLA_NET_0_74023);
    
    HIEFFPLA_INST_0_67878 : NOR3B
      port map(A => HIEFFPLA_NET_0_72743, B => 
        HIEFFPLA_NET_0_72895, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72781);
    
    HIEFFPLA_INST_0_56751 : AOI1C
      port map(A => HIEFFPLA_NET_0_75180, B => 
        HIEFFPLA_NET_0_75181, C => HIEFFPLA_NET_0_74754, Y => 
        HIEFFPLA_NET_0_75215);
    
    HIEFFPLA_INST_0_57654 : AOI1
      port map(A => \Science_0_exp_packet_0[34]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74979, Y => HIEFFPLA_NET_0_74980);
    
    HIEFFPLA_INST_0_57018 : AOI1D
      port map(A => HIEFFPLA_NET_0_74841, B => 
        HIEFFPLA_NET_0_74957, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75181);
    
    \Communications_0/UART_0/rx_clk_count[25]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75574, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75554, Q => 
        \Communications_0/UART_0/rx_clk_count[25]_net_1\);
    
    HIEFFPLA_INST_0_62064 : AND3C
      port map(A => HIEFFPLA_NET_0_74058, B => 
        HIEFFPLA_NET_0_74053, C => HIEFFPLA_NET_0_74048, Y => 
        HIEFFPLA_NET_0_74059);
    
    HIEFFPLA_INST_0_69233 : NOR3B
      port map(A => HIEFFPLA_NET_0_72454, B => 
        HIEFFPLA_NET_0_72488, C => HIEFFPLA_NET_0_72551, Y => 
        HIEFFPLA_NET_0_72442);
    
    \General_Controller_0/sweep_table_sweep_cnt[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74132, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[6]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/num_bytes_1[0]\ : 
        DFN1
      port map(D => HIEFFPLA_NET_0_72967, CLK => CLKINT_0_Y_0, Q
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[0]\);
    
    HIEFFPLA_INST_0_69003 : OR3B
      port map(A => HIEFFPLA_NET_0_72504, B => 
        HIEFFPLA_NET_0_72500, C => HIEFFPLA_NET_0_72487, Y => 
        HIEFFPLA_NET_0_72501);
    
    \General_Controller_0/en_data_saving\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74317, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74316, Q => 
        General_Controller_0_en_data_saving);
    
    HIEFFPLA_INST_0_57364 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_74854, Y => HIEFFPLA_NET_0_75066);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[12]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[12]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[12]\);
    
    HIEFFPLA_INST_0_60901 : OR3B
      port map(A => 
        \General_Controller_0/constant_bias_probe_id[0]_net_1\, B
         => HIEFFPLA_NET_0_74322, C => 
        \General_Controller_0/un10_uc_tx_rdy_i[1]\, Y => 
        HIEFFPLA_NET_0_74324);
    
    HIEFFPLA_INST_0_66644 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        C => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73075);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[3]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72263, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[3]_net_1\);
    
    \Science_0/ADC_READ_0/g4i[1]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73248, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73421, Q => 
        \Science_0/ADC_READ_0_G4[1]\);
    
    HIEFFPLA_INST_0_67162 : OR3B
      port map(A => HIEFFPLA_NET_0_72950, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[6]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72948);
    
    HIEFFPLA_INST_0_63698 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[3]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_nof_steps[3]_net_1\, S
         => \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73726);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_2[10]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74767, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\);
    
    HIEFFPLA_INST_0_60354 : MX2
      port map(A => \Sensors_0_acc_z[6]\, B => 
        \Sensors_0_acc_z[10]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74428);
    
    HIEFFPLA_INST_0_61627 : MX2
      port map(A => \SweepTable_0_RD[0]\, B => 
        \SweepTable_1_RD[0]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74170);
    
    HIEFFPLA_INST_0_61388 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[41]\, B => 
        \Timekeeper_0_milliseconds[1]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74205);
    
    HIEFFPLA_INST_0_71067 : AO1A
      port map(A => Communications_0_ext_tx_rdy, B => 
        HIEFFPLA_NET_0_71982, C => HIEFFPLA_NET_0_74605, Y => 
        HIEFFPLA_NET_0_74606);
    
    HIEFFPLA_INST_0_68025 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72751);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[20]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[20]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[20]\);
    
    \Science_0/SET_LP_GAIN_0/state[3]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73158, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/state_i_0[3]\);
    
    HIEFFPLA_INST_0_70508 : XOR2
      port map(A => HIEFFPLA_NET_0_72126, B => 
        \Timekeeper_0_milliseconds[21]\, Y => 
        HIEFFPLA_NET_0_72103);
    
    HIEFFPLA_INST_0_69044 : NAND2B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        Y => HIEFFPLA_NET_0_72487);
    
    HIEFFPLA_INST_0_57917 : AO1B
      port map(A => \Sensors_0_mag_time[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74905, Y => HIEFFPLA_NET_0_74906);
    
    \Communications_0/UART_0/tx_clk_count[6]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75520, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_clk_count_i_0[6]\);
    
    HIEFFPLA_INST_0_65492 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt2up[1]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2up[0]_net_1\, C => 
        HIEFFPLA_NET_0_73366, Y => HIEFFPLA_NET_0_73363);
    
    HIEFFPLA_INST_0_68143 : AO1
      port map(A => HIEFFPLA_NET_0_72747, B => 
        HIEFFPLA_NET_0_72762, C => HIEFFPLA_NET_0_72906, Y => 
        HIEFFPLA_NET_0_72724);
    
    HIEFFPLA_INST_0_67557 : OR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, B
         => HIEFFPLA_NET_0_72929, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72852);
    
    \Science_0/ADC_READ_0/exp_packet_1[22]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[6]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[22]\);
    
    HIEFFPLA_INST_0_65987 : NAND3
      port map(A => \Science_0/ADC_READ_0_G4[0]\, B => 
        \Science_0/ADC_READ_0/cnt4up[4]_net_1\, C => 
        HIEFFPLA_NET_0_73276, Y => HIEFFPLA_NET_0_73246);
    
    \FMC_DA_pad[3]/U0/U1\ : IOTRI_OB_EB
      port map(D => \FMC_DA_c[3]\, E => \VCC\, DOUT => 
        \FMC_DA_pad[3]/U0/NET1\, EOUT => \FMC_DA_pad[3]/U0/NET2\);
    
    \General_Controller_0/flight_state[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74290, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/flight_state[2]_net_1\);
    
    HIEFFPLA_INST_0_63860 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[6]_net_1\, B
         => 
        \General_Controller_0/sweep_table_sample_skip[6]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73699);
    
    \Science_0/ADC_READ_0/exp_packet_1[75]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[19]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[75]\);
    
    HIEFFPLA_INST_0_62969 : NAND3B
      port map(A => HIEFFPLA_NET_0_73785, B => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, C => 
        HIEFFPLA_NET_0_73987, Y => HIEFFPLA_NET_0_73855);
    
    \Science_0/ADC_READ_0/cnt3dn[1]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73346, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3dn[1]_net_1\);
    
    \Science_0/ADC_READ_0/chan7_data[11]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[17]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[11]\);
    
    HIEFFPLA_INST_0_58879 : AND3C
      port map(A => HIEFFPLA_NET_0_74697, B => 
        HIEFFPLA_NET_0_74650, C => HIEFFPLA_NET_0_74695, Y => 
        HIEFFPLA_NET_0_74667);
    
    HIEFFPLA_INST_0_64407 : MX2
      port map(A => HIEFFPLA_NET_0_73709, B => 
        HIEFFPLA_NET_0_73701, S => HIEFFPLA_NET_0_73593, Y => 
        HIEFFPLA_NET_0_73629);
    
    HIEFFPLA_INST_0_56612 : MX2
      port map(A => HIEFFPLA_NET_0_75199, B => 
        HIEFFPLA_NET_0_75069, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75232);
    
    HIEFFPLA_INST_0_66193 : AO1B
      port map(A => \Science_0/SET_LP_GAIN_0/state[6]_net_1\, B
         => \Science_0/ADC_READ_0_G2[1]\, C => 
        HIEFFPLA_NET_0_73181, Y => HIEFFPLA_NET_0_73182);
    
    \ACCE_SDA_pad/U0/U1\ : IOBI_IB_OB_EB
      port map(D => 
        \Sensors_0.Accelerometer_0.I2C_Master_0.sda_1\, E => 
        sda_cl_1_RNIBFPP, YIN => \ACCE_SDA_pad/U0/NET3\, DOUT => 
        \ACCE_SDA_pad/U0/NET1\, EOUT => \ACCE_SDA_pad/U0/NET2\, Y
         => ACCE_SDA_in);
    
    HIEFFPLA_INST_0_58536 : XA1
      port map(A => HIEFFPLA_NET_0_74727, B => 
        \Eject_Signal_Debounce_0/ms_cnt[5]_net_1\, C => 
        HIEFFPLA_NET_0_74738, Y => HIEFFPLA_NET_0_74741);
    
    HIEFFPLA_INST_0_68504 : AND3C
      port map(A => HIEFFPLA_NET_0_72707, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[0]_net_1\, C => 
        HIEFFPLA_NET_0_72625, Y => HIEFFPLA_NET_0_72634);
    
    HIEFFPLA_INST_0_58543 : NAND3A
      port map(A => CLKINT_1_Y, B => 
        \Eject_Signal_Debounce_0/old_1kHz_i_0\, C => \m_time[7]\, 
        Y => HIEFFPLA_NET_0_74739);
    
    HIEFFPLA_INST_0_63704 : MX2
      port map(A => 
        \General_Controller_0/constant_bias_voltage_0[4]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_nof_steps[4]_net_1\, S
         => \General_Controller_0/uc_tx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73725);
    
    HIEFFPLA_INST_0_68862 : AO1A
      port map(A => HIEFFPLA_NET_0_72501, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[2]_net_1\, C
         => HIEFFPLA_NET_0_72536, Y => HIEFFPLA_NET_0_72537);
    
    HIEFFPLA_INST_0_64979 : OR3B
      port map(A => HIEFFPLA_NET_0_73499, B => 
        \Pressure_Signal_Debounce_0/ms_cnt[8]_net_1\, C => 
        HIEFFPLA_NET_0_73500, Y => HIEFFPLA_NET_0_73496);
    
    HIEFFPLA_INST_0_71118 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_71979, Y => HIEFFPLA_NET_0_75014);
    
    \Data_Saving_0/Packet_Saver_0/old_pressure_new_data\ : DFN0P1
      port map(D => \AFLSDF_INV_33\, CLK => CLKINT_0_Y_0, PRE => 
        CLKINT_1_Y, Q => 
        \Data_Saving_0/Packet_Saver_0/old_pressure_new_data_i_0\);
    
    HIEFFPLA_INST_0_58444 : OA1C
      port map(A => HIEFFPLA_NET_0_74767, B => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, C => 
        HIEFFPLA_NET_0_74764, Y => HIEFFPLA_NET_0_74765);
    
    HIEFFPLA_INST_0_68429 : MX2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[3]\, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[7]\, S => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72652);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73141, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\);
    
    HIEFFPLA_INST_0_59187 : NOR3B
      port map(A => \GS_Readout_0/state[6]_net_1\, B => 
        \GS_Readout_0/prevState[1]_net_1\, C => 
        Communications_0_ext_tx_rdy, Y => HIEFFPLA_NET_0_74593);
    
    HIEFFPLA_INST_0_59229 : NOR3B
      port map(A => \GS_Readout_0/prevState[5]_net_1\, B => 
        HIEFFPLA_NET_0_74718, C => 
        \GS_Readout_0/prevState[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74584);
    
    HIEFFPLA_INST_0_57282 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[52]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_75098);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_RGRY[3]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75302, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[3]\\\\\);
    
    \Communications_0/UART_0/tx_count[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75505, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75503, Q => 
        \Communications_0/UART_0/tx_count[2]_net_1\);
    
    HIEFFPLA_INST_0_63496 : MX2
      port map(A => HIEFFPLA_NET_0_73682, B => 
        HIEFFPLA_NET_0_73674, S => HIEFFPLA_NET_0_73621, Y => 
        HIEFFPLA_NET_0_73757);
    
    HIEFFPLA_INST_0_61924 : AND3
      port map(A => HIEFFPLA_NET_0_74113, B => 
        HIEFFPLA_NET_0_74091, C => HIEFFPLA_NET_0_74079, Y => 
        HIEFFPLA_NET_0_74097);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/data_out[6]\ : 
        DFN0E1C1
      port map(D => ACCE_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73117, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[6]\);
    
    \Science_0/ADC_READ_0/chan1_data[11]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[17]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[11]\);
    
    HIEFFPLA_INST_0_58959 : NOR3B
      port map(A => HIEFFPLA_NET_0_74564, B => 
        \GS_Readout_0/state[2]_net_1\, C => HIEFFPLA_NET_0_74725, 
        Y => HIEFFPLA_NET_0_74649);
    
    HIEFFPLA_INST_0_63000 : AOI1B
      port map(A => HIEFFPLA_NET_0_73887, B => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, C => 
        HIEFFPLA_NET_0_74037, Y => HIEFFPLA_NET_0_73850);
    
    HIEFFPLA_INST_0_70503 : XOR2
      port map(A => HIEFFPLA_NET_0_72123, B => 
        \Timekeeper_0_milliseconds[19]\, Y => 
        HIEFFPLA_NET_0_72106);
    
    \Timing_0/m_count[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72080, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_count[0]_net_1\);
    
    \Science_0/ADC_READ_0/data_a[3]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[2]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[3]_net_1\);
    
    HIEFFPLA_INST_0_57270 : AND2
      port map(A => \Sensors_0_gyro_time[14]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75101);
    
    HIEFFPLA_INST_0_54983 : XO1
      port map(A => \Communications_0/UART_0_recv[1]\, B => 
        \General_Controller_0_unit_id[1]\, C => 
        HIEFFPLA_NET_0_75620, Y => HIEFFPLA_NET_0_75621);
    
    HIEFFPLA_INST_0_56514 : AND2
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, B
         => HIEFFPLA_NET_0_75349, Y => HIEFFPLA_NET_0_75257);
    
    HIEFFPLA_INST_0_67554 : OR2A
      port map(A => HIEFFPLA_NET_0_72741, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, Y
         => HIEFFPLA_NET_0_72853);
    
    HIEFFPLA_INST_0_65618 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt4dn[2]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt4dn[0]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt4dn[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73329);
    
    \Eject_Signal_Debounce_0/ms_cnt[3]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74743, CLK => CLKINT_0_Y_0, Q
         => \Eject_Signal_Debounce_0/ms_cnt[3]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72728, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\);
    
    HIEFFPLA_INST_0_67306 : AND2B
      port map(A => HIEFFPLA_NET_0_72935, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72911);
    
    HIEFFPLA_INST_0_56069 : XA1A
      port map(A => HIEFFPLA_NET_0_75328, B => 
        HIEFFPLA_NET_0_75258, C => HIEFFPLA_NET_0_75355, Y => 
        HIEFFPLA_NET_0_75356);
    
    HIEFFPLA_INST_0_64454 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state[4]_net_1\, 
        B => HIEFFPLA_NET_0_74037, C => 
        \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73623);
    
    HIEFFPLA_INST_0_66068 : AX1D
      port map(A => \Science_0/DAC_SET_0/state[3]_net_1\, B => 
        \Science_0/DAC_SET_0/state[1]_net_1\, C => 
        \Science_0/DAC_SET_0/cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73219);
    
    HIEFFPLA_INST_0_57292 : AND2
      port map(A => \Sensors_0_mag_y[8]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        Y => HIEFFPLA_NET_0_75088);
    
    HIEFFPLA_INST_0_66941 : AO1D
      port map(A => HIEFFPLA_NET_0_72738, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        C => HIEFFPLA_NET_0_72929, Y => HIEFFPLA_NET_0_73000);
    
    HIEFFPLA_INST_0_62474 : NOR3B
      port map(A => \General_Controller_0/uc_rx_state[2]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[4]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73975);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[2]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72279, Q => 
        \Sensors_0_pressure_temp_raw[2]\);
    
    \General_Controller_0/sweep_table_write_value[0]\ : DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[0]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[0]_net_1\);
    
    \General_Controller_0/st_wdata[14]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[14]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[14]\);
    
    \General_Controller_0/status_bits_1[60]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74186, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[60]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[55]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/chan[1]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[55]\);
    
    \Science_0/ADC_READ_0/chan6_data[11]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[17]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[11]\);
    
    HIEFFPLA_INST_0_62221 : NOR3A
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state[4]_net_1\, C => 
        \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74026);
    
    HIEFFPLA_INST_0_61743 : AND3
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[9]_net_1\, B
         => HIEFFPLA_NET_0_74146, C => 
        \General_Controller_0/sweep_table_sweep_cnt[10]_net_1\, Y
         => HIEFFPLA_NET_0_74149);
    
    HIEFFPLA_INST_0_60872 : OR3A
      port map(A => \General_Controller_0/command[0]_net_1\, B
         => HIEFFPLA_NET_0_74329, C => HIEFFPLA_NET_0_74335, Y
         => HIEFFPLA_NET_0_74334);
    
    HIEFFPLA_INST_0_66802 : AO1A
      port map(A => HIEFFPLA_NET_0_73101, B => 
        HIEFFPLA_NET_0_73059, C => HIEFFPLA_NET_0_73031, Y => 
        HIEFFPLA_NET_0_73032);
    
    \Sensors_0/Gyro_0/I2C_Master_0/write_done\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72629, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72571, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_write_done\);
    
    \Science_0/ADC_READ_0/cnt[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73285, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73242, Q => 
        \Science_0/ADC_READ_0/cnt[5]_net_1\);
    
    HIEFFPLA_INST_0_57129 : AO1
      port map(A => \Sensors_0_acc_time[13]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_75102, Y => HIEFFPLA_NET_0_75164);
    
    \Science_0/ADC_READ_0/chan6_data[7]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[7]\);
    
    \Science_0/ADC_READ_0/chan0_data[7]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[7]\);
    
    HIEFFPLA_INST_0_65748 : AND2A
      port map(A => HIEFFPLA_NET_0_73241, B => 
        HIEFFPLA_NET_0_73289, Y => HIEFFPLA_NET_0_73290);
    
    HIEFFPLA_INST_0_56527 : XNOR2
      port map(A => 
        \Data_Saving_0/Interrupt_Generator_0/counter[0]_net_1\, B
         => CLKINT_1_Y, Y => HIEFFPLA_NET_0_75253);
    
    \General_Controller_0/sweep_table_read_value[15]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74164, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[15]_net_1\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[0]\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_73130, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73041, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[0]_net_1\);
    
    HIEFFPLA_INST_0_70208 : AND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[5]_net_1\, 
        B => \Sensors_0/Pressure_Sensor_0/state[8]\, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72196);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[9]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72777, Q => 
        \Sensors_0_acc_y[9]\);
    
    HIEFFPLA_INST_0_68291 : MX2A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[0]_net_1\, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_num_bytes[0]\, S
         => \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_72688);
    
    HIEFFPLA_INST_0_61730 : XA1B
      port map(A => HIEFFPLA_NET_0_73539, B => 
        \General_Controller_0/sweep_table_read_wait[30]_net_1\, C
         => HIEFFPLA_NET_0_73977, Y => HIEFFPLA_NET_0_74152);
    
    HIEFFPLA_INST_0_65218 : AND3
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[1]_net_1\, 
        B => \Pressure_Signal_Debounce_0/ms_cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_73478, Y => HIEFFPLA_NET_0_73443);
    
    HIEFFPLA_INST_0_60288 : NOR3B
      port map(A => HIEFFPLA_NET_0_74490, B => 
        HIEFFPLA_NET_0_74450, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74436);
    
    \General_Controller_0/constant_bias_voltage_0[7]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[7]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[7]_net_1\);
    
    HIEFFPLA_INST_0_55353 : AND2
      port map(A => \Communications_0/UART_0/tx_clk_count_i_0[2]\, 
        B => \Communications_0/UART_0/tx_clk_count_i_0[3]\, Y => 
        HIEFFPLA_NET_0_75532);
    
    HIEFFPLA_INST_0_65416 : OR3A
      port map(A => HIEFFPLA_NET_0_73277, B => 
        HIEFFPLA_NET_0_73383, C => HIEFFPLA_NET_0_73385, Y => 
        HIEFFPLA_NET_0_73382);
    
    \Science_0/ADC_READ_0/cnt2dn[4]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73372, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2dn[4]_net_1\);
    
    HIEFFPLA_INST_0_69157 : NOR3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\, 
        B => HIEFFPLA_NET_0_72544, C => 
        \Sensors_0/Gyro_0/I2C_Master_0_write_done\, Y => 
        HIEFFPLA_NET_0_72458);
    
    HIEFFPLA_INST_0_63824 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[0]_net_1\, B
         => 
        \General_Controller_0/sweep_table_sample_skip[0]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73705);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/write_done\ : 
        DFN0E1C1
      port map(D => HIEFFPLA_NET_0_73050, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73009, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\);
    
    HIEFFPLA_INST_0_62382 : AND3B
      port map(A => HIEFFPLA_NET_0_74007, B => 
        HIEFFPLA_NET_0_74005, C => HIEFFPLA_NET_0_73783, Y => 
        HIEFFPLA_NET_0_73993);
    
    HIEFFPLA_INST_0_58513 : XA1
      port map(A => \Eject_Signal_Debounce_0/ms_cnt[1]_net_1\, B
         => HIEFFPLA_NET_0_74733, C => HIEFFPLA_NET_0_74738, Y
         => HIEFFPLA_NET_0_74745);
    
    HIEFFPLA_INST_0_57155 : AND2
      port map(A => \Sensors_0_pressure_time[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, Y
         => HIEFFPLA_NET_0_75150);
    
    HIEFFPLA_INST_0_58953 : NOR3B
      port map(A => HIEFFPLA_NET_0_74368, B => 
        HIEFFPLA_NET_0_74647, C => HIEFFPLA_NET_0_74360, Y => 
        HIEFFPLA_NET_0_74650);
    
    \General_Controller_0/sweep_table_samples_per_step[5]\ : 
        DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[5]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[5]_net_1\);
    
    \Pressure_Signal_Debounce_0/ms_cnt[0]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73495, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[0]_net_1\);
    
    HIEFFPLA_INST_0_58998 : NOR2A
      port map(A => \GS_Readout_0/state[3]_net_1\, B => 
        HIEFFPLA_NET_0_74372, Y => HIEFFPLA_NET_0_74641);
    
    HIEFFPLA_INST_0_62162 : AND2B
      port map(A => HIEFFPLA_NET_0_73933, B => 
        HIEFFPLA_NET_0_73977, Y => HIEFFPLA_NET_0_74039);
    
    HIEFFPLA_INST_0_67858 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72786);
    
    HIEFFPLA_INST_0_66521 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]_net_1\, 
        B => ACCE_SCL_c, C => HIEFFPLA_NET_0_73145, Y => 
        HIEFFPLA_NET_0_73103);
    
    HIEFFPLA_INST_0_57509 : AO1B
      port map(A => \Sensors_0_mag_z[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75024, Y => HIEFFPLA_NET_0_75025);
    
    HIEFFPLA_INST_0_69558 : AO1A
      port map(A => HIEFFPLA_NET_0_72429, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[1]\, 
        C => HIEFFPLA_NET_0_72374, Y => HIEFFPLA_NET_0_72365);
    
    HIEFFPLA_INST_0_62095 : NOR3B
      port map(A => HIEFFPLA_NET_0_73890, B => 
        HIEFFPLA_NET_0_74018, C => 
        \General_Controller_0/uc_rx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74053);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[17]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[17]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[17]\);
    
    HIEFFPLA_INST_0_65998 : NOR2A
      port map(A => \Science_0/ADC_READ_0/newflag_net_1\, B => 
        HIEFFPLA_NET_0_73414, Y => HIEFFPLA_NET_0_73244);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[10]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[10]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[10]\);
    
    HIEFFPLA_INST_0_57380 : AO1
      port map(A => \Science_0_exp_packet_0[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74852, Y => HIEFFPLA_NET_0_75062);
    
    \Communications_0/UART_1/rx_clk_count[27]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75460, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75443, Q => 
        \Communications_0/UART_1/rx_clk_count[27]_net_1\);
    
    HIEFFPLA_INST_0_57827 : AO1B
      port map(A => \Sensors_0_mag_time[18]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74932, Y => HIEFFPLA_NET_0_74933);
    
    \General_Controller_0/sweep_table_samples_per_step[13]\ : 
        DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[13]_net_1\);
    
    HIEFFPLA_INST_0_70197 : OA1A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        B => HIEFFPLA_NET_0_72187, C => HIEFFPLA_NET_0_72186, Y
         => HIEFFPLA_NET_0_72197);
    
    HIEFFPLA_INST_0_61675 : MX2
      port map(A => \SweepTable_0_RD[2]\, B => 
        \SweepTable_1_RD[2]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74162);
    
    \Data_Saving_0/Packet_Saver_0/gyro_flag\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_74774, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => 
        General_Controller_0_en_data_saving, Q => 
        \Data_Saving_0/Packet_Saver_0/gyro_flag_net_1\);
    
    HIEFFPLA_INST_0_64114 : OR2A
      port map(A => HIEFFPLA_NET_0_73579, B => 
        \General_Controller_0/constant_bias_voltage_0[13]_net_1\, 
        Y => HIEFFPLA_NET_0_73667);
    
    \General_Controller_0/sweep_table_read_value[12]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74167, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[12]_net_1\);
    
    HIEFFPLA_INST_0_70585 : AX1C
      port map(A => HIEFFPLA_NET_0_72032, B => 
        HIEFFPLA_NET_0_72030, C => \Timing_0/m_count[6]_net_1\, Y
         => HIEFFPLA_NET_0_72072);
    
    HIEFFPLA_INST_0_70217 : AO1A
      port map(A => HIEFFPLA_NET_0_72273, B => 
        HIEFFPLA_NET_0_72184, C => HIEFFPLA_NET_0_72234, Y => 
        HIEFFPLA_NET_0_72193);
    
    HIEFFPLA_INST_0_67800 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, B
         => HIEFFPLA_NET_0_72739, C => HIEFFPLA_NET_0_72799, Y
         => HIEFFPLA_NET_0_72798);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_time[15]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[15]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72923, Q => 
        \Sensors_0_mag_time[15]\);
    
    HIEFFPLA_INST_0_61739 : AND3
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[3]_net_1\, B
         => HIEFFPLA_NET_0_74148, C => 
        \General_Controller_0/sweep_table_sweep_cnt[4]_net_1\, Y
         => HIEFFPLA_NET_0_74150);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[11]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72807, Q => 
        \Sensors_0_mag_z[11]\);
    
    HIEFFPLA_INST_0_64857 : MX2
      port map(A => HIEFFPLA_NET_0_73527, B => 
        HIEFFPLA_NET_0_73582, S => Communications_0_uc_tx_rdy, Y
         => HIEFFPLA_NET_0_73523);
    
    HIEFFPLA_INST_0_57216 : AND2
      port map(A => \Sensors_0_acc_time[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, Y
         => HIEFFPLA_NET_0_75125);
    
    HIEFFPLA_INST_0_55431 : AX1B
      port map(A => HIEFFPLA_NET_0_75501, B => 
        HIEFFPLA_NET_0_75533, C => 
        \Communications_0/UART_0/tx_clk_count_i_0[2]\, Y => 
        HIEFFPLA_NET_0_75515);
    
    HIEFFPLA_INST_0_70259 : AO1D
      port map(A => HIEFFPLA_NET_0_72308, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        C => HIEFFPLA_NET_0_72302, Y => HIEFFPLA_NET_0_72185);
    
    HIEFFPLA_INST_0_68619 : AND3C
      port map(A => HIEFFPLA_NET_0_72598, B => 
        HIEFFPLA_NET_0_72595, C => HIEFFPLA_NET_0_72593, Y => 
        HIEFFPLA_NET_0_72604);
    
    HIEFFPLA_INST_0_60929 : MX2A
      port map(A => General_Controller_0_en_data_saving, B => 
        \General_Controller_0/flight_state[2]_net_1\, S => 
        HIEFFPLA_NET_0_74337, Y => HIEFFPLA_NET_0_74317);
    
    \General_Controller_0/sweep_table_read_value[0]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74170, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[0]_net_1\);
    
    HIEFFPLA_INST_0_59103 : AO1A
      port map(A => HIEFFPLA_NET_0_74382, B => 
        \GS_Readout_0/state[2]_net_1\, C => HIEFFPLA_NET_0_74611, 
        Y => HIEFFPLA_NET_0_74612);
    
    \Timekeeper_0/milliseconds[13]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72112, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[13]\);
    
    \Science_0/ADC_READ_0/data_b[4]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[3]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[4]_net_1\);
    
    HIEFFPLA_INST_0_61919 : AND3B
      port map(A => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        B => \General_Controller_0/uc_rx_byte[3]_net_1\, C => 
        HIEFFPLA_NET_0_74098, Y => HIEFFPLA_NET_0_74099);
    
    \General_Controller_0/status_bits_1[53]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74193, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[53]\);
    
    HIEFFPLA_INST_0_65555 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt3dn[3]_net_1\, B => 
        HIEFFPLA_NET_0_73348, C => HIEFFPLA_NET_0_73349, Y => 
        HIEFFPLA_NET_0_73344);
    
    HIEFFPLA_INST_0_64108 : OR2A
      port map(A => HIEFFPLA_NET_0_73579, B => 
        \General_Controller_0/constant_bias_voltage_0[8]_net_1\, 
        Y => HIEFFPLA_NET_0_73670);
    
    \Science_0/ADC_READ_0/cnt4up[1]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73305, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4up[1]_net_1\);
    
    HIEFFPLA_INST_0_62733 : NAND2A
      port map(A => HIEFFPLA_NET_0_73904, B => 
        HIEFFPLA_NET_0_73934, Y => HIEFFPLA_NET_0_73919);
    
    HIEFFPLA_INST_0_70511 : AX1C
      port map(A => HIEFFPLA_NET_0_72126, B => 
        \Timekeeper_0_milliseconds[21]\, C => 
        \Timekeeper_0_milliseconds[22]\, Y => 
        HIEFFPLA_NET_0_72102);
    
    HIEFFPLA_INST_0_69416 : NAND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72394);
    
    HIEFFPLA_INST_0_58318 : AO1
      port map(A => \Sensors_0_mag_y[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75084, Y => HIEFFPLA_NET_0_74803);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72213, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\);
    
    HIEFFPLA_INST_0_61356 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[0]\, B => 
        \General_Controller_0/mission_mode_net_1\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74209);
    
    \UC_I2C4_SDA_pad/U0/U0\ : IOPAD_BI
      port map(D => \UC_I2C4_SDA_pad/U0/NET1\, E => 
        \UC_I2C4_SDA_pad/U0/NET2\, Y => \UC_I2C4_SDA_pad/U0/NET3\, 
        PAD => UC_I2C4_SDA);
    
    \L2WR_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => L2WR_c, E => \VCC\, DOUT => 
        \L2WR_pad/U0/NET1\, EOUT => \L2WR_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_70749 : AX1C
      port map(A => HIEFFPLA_NET_0_72026, B => 
        \Timing_0/s_count[1]_net_1\, C => 
        \Timing_0/s_count[2]_net_1\, Y => HIEFFPLA_NET_0_72023);
    
    \General_Controller_0/st_wdata[8]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[8]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[8]\);
    
    HIEFFPLA_INST_0_71017 : OA1A
      port map(A => \General_Controller_0/uc_tx_state[4]_net_1\, 
        B => \General_Controller_0/uc_tx_substate[1]_net_1\, C
         => HIEFFPLA_NET_0_73592, Y => HIEFFPLA_NET_0_71987);
    
    HIEFFPLA_INST_0_64815 : AND3
      port map(A => HIEFFPLA_NET_0_73780, B => 
        HIEFFPLA_NET_0_74013, C => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73535);
    
    HIEFFPLA_INST_0_63214 : NOR3A
      port map(A => HIEFFPLA_NET_0_73907, B => 
        HIEFFPLA_NET_0_73811, C => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73805);
    
    \ARST_pad/U0/U0\ : IOPAD_TRI
      port map(D => \ARST_pad/U0/NET1\, E => \ARST_pad/U0/NET2\, 
        PAD => ARST);
    
    HIEFFPLA_INST_0_57963 : AO1
      port map(A => \Science_0_exp_packet_0[71]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_74789, Y => HIEFFPLA_NET_0_74892);
    
    \Science_0/SET_LP_GAIN_0/old_G4[1]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73162, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/old_G4[1]_net_1\);
    
    HIEFFPLA_INST_0_57228 : AND2
      port map(A => \Sensors_0_pressure_time[16]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75120);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_x[0]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72801, Q => 
        \Sensors_0_acc_x[0]\);
    
    HIEFFPLA_INST_0_64954 : AX1C
      port map(A => \I2C_PassThrough_0/cnt[0]_net_1\, B => 
        HIEFFPLA_NET_0_73514, C => 
        \I2C_PassThrough_0/cnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73504);
    
    HIEFFPLA_INST_0_59403 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[42]\, B => 
        \Data_Hub_Packets_0_status_packet[46]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74559);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[10]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72484, Q => 
        \Sensors_0_gyro_y[10]\);
    
    \FMC_CLK_pad/U0/U1\ : IOIN_IB
      port map(YIN => \FMC_CLK_pad/U0/NET1\, Y => FMC_CLK_c);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73035, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\);
    
    \I2C_PassThrough_0/state[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73511, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \I2C_PassThrough_0.state[2]\);
    
    AFLSDF_INV_15 : INV
      port map(A => CLKINT_1_Y, Y => \AFLSDF_INV_15\);
    
    HIEFFPLA_INST_0_69053 : NOR3B
      port map(A => HIEFFPLA_NET_0_72483, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[6]_net_1\, 
        C => HIEFFPLA_NET_0_72548, Y => HIEFFPLA_NET_0_72484);
    
    HIEFFPLA_INST_0_62974 : NOR3A
      port map(A => HIEFFPLA_NET_0_73885, B => 
        HIEFFPLA_NET_0_73987, C => 
        \General_Controller_0/uc_rx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73854);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_1[12]\ : DFN0E0P1
      port map(D => HIEFFPLA_NET_0_75241, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\);
    
    \General_Controller_0/uc_tx_nextstate[7]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73931, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73857, Q => 
        \General_Controller_0/uc_tx_nextstate[7]_net_1\);
    
    \Science_0/ADC_READ_0/chan7_data[7]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[13]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[7]\);
    
    HIEFFPLA_INST_0_57250 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[57]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_75113);
    
    HIEFFPLA_INST_0_65138 : AO1A
      port map(A => \Sensors_0_pressure_raw[1]\, B => 
        HIEFFPLA_NET_0_73469, C => HIEFFPLA_NET_0_73457, Y => 
        HIEFFPLA_NET_0_73461);
    
    HIEFFPLA_INST_0_56857 : MX2
      port map(A => HIEFFPLA_NET_0_75008, B => 
        HIEFFPLA_NET_0_74934, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75203);
    
    HIEFFPLA_INST_0_59306 : MX2
      port map(A => HIEFFPLA_NET_0_74342, B => 
        HIEFFPLA_NET_0_74487, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74571);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[7]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72503, Q => 
        \Sensors_0_gyro_x[7]\);
    
    \Pressure_Signal_Debounce_0/ms_cnt[3]\ : DFN1
      port map(D => HIEFFPLA_NET_0_73492, CLK => \m_time[7]\, Q
         => \Pressure_Signal_Debounce_0/ms_cnt[3]_net_1\);
    
    HIEFFPLA_INST_0_70012 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_72228, C => HIEFFPLA_NET_0_72243, Y
         => HIEFFPLA_NET_0_72247);
    
    HIEFFPLA_INST_0_55420 : AOI1D
      port map(A => \Communications_0/UART_0/tx_clk_count_i_0[7]\, 
        B => HIEFFPLA_NET_0_75535, C => 
        \Communications_0/UART_0/tx_clk_count_i_0[8]\, Y => 
        HIEFFPLA_NET_0_75517);
    
    HIEFFPLA_INST_0_61790 : XOR2
      port map(A => HIEFFPLA_NET_0_74145, B => 
        \General_Controller_0/sweep_table_sweep_cnt[7]_net_1\, Y
         => HIEFFPLA_NET_0_74131);
    
    HIEFFPLA_INST_0_67927 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72771);
    
    HIEFFPLA_INST_0_63662 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[13]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_samples_per_point[13]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73732);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[3]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[3]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[3]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[17]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[17]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[17]\);
    
    HIEFFPLA_INST_0_62742 : XA1
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_73860, Y => HIEFFPLA_NET_0_73917);
    
    HIEFFPLA_INST_0_60039 : MX2
      port map(A => HIEFFPLA_NET_0_74515, B => 
        HIEFFPLA_NET_0_74491, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74470);
    
    \Communications_0/FFU_Command_Checker_0/command_out[1]\ : 
        DFN1E1C1
      port map(D => \Communications_0/UART_0_recv[1]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75625, Q => \Communications_0_ext_recv[1]\);
    
    HIEFFPLA_INST_0_69084 : OR3B
      port map(A => HIEFFPLA_NET_0_72504, B => 
        HIEFFPLA_NET_0_72473, C => HIEFFPLA_NET_0_72487, Y => 
        HIEFFPLA_NET_0_72474);
    
    HIEFFPLA_INST_0_61230 : NAND3C
      port map(A => \General_Controller_0/state_seconds[9]_net_1\, 
        B => \General_Controller_0/state_seconds[18]_net_1\, C
         => \General_Controller_0/state_seconds[11]_net_1\, Y => 
        HIEFFPLA_NET_0_74242);
    
    HIEFFPLA_INST_0_57211 : AND2
      port map(A => \Sensors_0_gyro_y[14]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75128);
    
    HIEFFPLA_INST_0_67821 : AO1
      port map(A => HIEFFPLA_NET_0_72759, B => 
        HIEFFPLA_NET_0_72881, C => HIEFFPLA_NET_0_72788, Y => 
        HIEFFPLA_NET_0_72794);
    
    HIEFFPLA_INST_0_59124 : AO1A
      port map(A => HIEFFPLA_NET_0_74382, B => 
        \GS_Readout_0/state[4]_net_1\, C => HIEFFPLA_NET_0_74606, 
        Y => HIEFFPLA_NET_0_74607);
    
    HIEFFPLA_INST_0_69327 : NAND2B
      port map(A => HIEFFPLA_NET_0_72415, B => 
        HIEFFPLA_NET_0_72319, Y => HIEFFPLA_NET_0_72417);
    
    \I2C_PassThrough_0/state[3]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73510, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \I2C_PassThrough_0.state[3]\);
    
    HIEFFPLA_INST_0_69605 : NAND3C
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[7]_net_1\, 
        B => HIEFFPLA_NET_0_72341, C => HIEFFPLA_NET_0_72422, Y
         => HIEFFPLA_NET_0_72352);
    
    \Communications_0/UART_0/recv[6]\ : DFN1E1C1
      port map(D => \Communications_0/UART_0/rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75551, Q => 
        \Communications_0/UART_0_recv[6]\);
    
    \UC_RESET_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => \GND\, E => \GND\, DOUT => 
        \UC_RESET_pad/U0/NET1\, EOUT => \UC_RESET_pad/U0/NET2\);
    
    HIEFFPLA_INST_0_63269 : AND2B
      port map(A => HIEFFPLA_NET_0_73917, B => 
        HIEFFPLA_NET_0_73812, Y => HIEFFPLA_NET_0_73794);
    
    \Science_0/ADC_READ_0/cnt4dn[6]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73312, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4dn[6]_net_1\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72694, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\);
    
    HIEFFPLA_INST_0_67261 : AO1
      port map(A => HIEFFPLA_NET_0_72805, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        Y => HIEFFPLA_NET_0_72924);
    
    \General_Controller_0/st_raddr[6]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73979, Q => 
        \General_Controller_0_st_raddr_1[6]\);
    
    \Science_0/ADC_READ_0/chan2_data[0]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[0]\);
    
    HIEFFPLA_INST_0_62368 : NOR3B
      port map(A => HIEFFPLA_NET_0_73995, B => 
        HIEFFPLA_NET_0_74113, C => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73996);
    
    HIEFFPLA_INST_0_68836 : NAND2B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, B
         => HIEFFPLA_NET_0_72540, Y => HIEFFPLA_NET_0_72544);
    
    HIEFFPLA_INST_0_69807 : XA1
      port map(A => HIEFFPLA_NET_0_72306, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[2]_net_1\, 
        C => HIEFFPLA_NET_0_72236, Y => HIEFFPLA_NET_0_72298);
    
    \Science_0/SET_LP_GAIN_0/old_G4[0]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73164, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/old_G4[0]_net_1\);
    
    HIEFFPLA_INST_0_69380 : XOR2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72403);
    
    HIEFFPLA_INST_0_70539 : AX1C
      port map(A => \Timing_0/f_time[0]_net_1\, B => 
        \Timing_0/f_time[1]_net_1\, C => 
        \Timing_0/f_time[2]_net_1\, Y => HIEFFPLA_NET_0_72088);
    
    HIEFFPLA_INST_0_58342 : AO1
      port map(A => \Sensors_0_mag_x[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75094, Y => HIEFFPLA_NET_0_74797);
    
    \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]\ : DFN0E0
      port map(D => HIEFFPLA_NET_0_72667, CLK => 
        ClockDivs_0_clk_800kHz, E => HIEFFPLA_NET_0_72617, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[1]_net_1\);
    
    HIEFFPLA_INST_0_66214 : MX2
      port map(A => \Science_0/SET_LP_GAIN_0/old_G1[1]_net_1\, B
         => \Science_0/ADC_READ_0_G1[1]\, S => 
        \Science_0/SET_LP_GAIN_0/state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73176);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_17\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[8]\\\\\, CLK => 
        CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_17_Q\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_WADDR[1]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75294, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[1]\\\\\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[4]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[4]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[4]\);
    
    \General_Controller_0/st_wen0\ : DFI1E1C1
      port map(D => HIEFFPLA_NET_0_74179, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_74177, CLR => CLKINT_1_Y, QN => 
        \SweepTable_0.WEAP\);
    
    HIEFFPLA_INST_0_70695 : XOR2
      port map(A => \Timing_0/s_time[8]_net_1\, B => 
        HIEFFPLA_NET_0_72037, Y => HIEFFPLA_NET_0_72041);
    
    HIEFFPLA_INST_0_65875 : AO1A
      port map(A => HIEFFPLA_NET_0_73263, B => 
        HIEFFPLA_NET_0_73261, C => HIEFFPLA_NET_0_73265, Y => 
        HIEFFPLA_NET_0_73266);
    
    HIEFFPLA_INST_0_56391 : AX1D
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, B
         => HIEFFPLA_NET_0_75351, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\, Y
         => HIEFFPLA_NET_0_75292);
    
    HIEFFPLA_INST_0_55009 : XO1
      port map(A => \Communications_0/UART_0_recv[7]\, B => 
        \General_Controller_0_unit_id[7]\, C => 
        HIEFFPLA_NET_0_75613, Y => HIEFFPLA_NET_0_75617);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[6]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72919, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[6]_net_1\);
    
    HIEFFPLA_INST_0_67890 : AO1
      port map(A => HIEFFPLA_NET_0_72802, B => 
        HIEFFPLA_NET_0_72929, C => HIEFFPLA_NET_0_72787, Y => 
        HIEFFPLA_NET_0_72779);
    
    \Timing_0/s_time[9]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72043, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \s_clks_net_0[24]\);
    
    HIEFFPLA_INST_0_58076 : AND2
      port map(A => \ch3_data_net_0[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_74862);
    
    HIEFFPLA_INST_0_69348 : AND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/next_state[2]_net_1\, 
        B => HIEFFPLA_NET_0_72410, Y => HIEFFPLA_NET_0_72412);
    
    HIEFFPLA_INST_0_69989 : NOR3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/isSetup_net_1\, 
        C => HIEFFPLA_NET_0_72245, Y => HIEFFPLA_NET_0_72251);
    
    HIEFFPLA_INST_0_69020 : AND2
      port map(A => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72496);
    
    HIEFFPLA_INST_0_66675 : AO1
      port map(A => HIEFFPLA_NET_0_73132, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        C => HIEFFPLA_NET_0_73142, Y => HIEFFPLA_NET_0_73068);
    
    \Science_0/ADC_READ_0/exp_packet_1[18]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_b[2]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[18]\);
    
    HIEFFPLA_INST_0_57376 : AO1
      port map(A => \Sensors_0_gyro_temp[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75062, Y => HIEFFPLA_NET_0_75063);
    
    \Science_0/ADC_RESET_0/ADCRESET\ : DFN1C1
      port map(D => \Science_0/ADC_RESET_0/state[1]_net_1\, CLK
         => \s_time[5]\, CLR => CLKINT_1_Y, Q => ARST_c);
    
    HIEFFPLA_INST_0_66713 : OR3A
      port map(A => HIEFFPLA_NET_0_73057, B => 
        HIEFFPLA_NET_0_73038, C => HIEFFPLA_NET_0_73062, Y => 
        HIEFFPLA_NET_0_73056);
    
    HIEFFPLA_INST_0_60122 : MX2
      port map(A => \Science_0_chan2_data[4]\, B => 
        \Science_0_chan2_data[8]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74458);
    
    HIEFFPLA_INST_0_67489 : NAND3C
      port map(A => HIEFFPLA_NET_0_72854, B => 
        HIEFFPLA_NET_0_72945, C => HIEFFPLA_NET_0_72834, Y => 
        HIEFFPLA_NET_0_72866);
    
    HIEFFPLA_INST_0_61850 : NAND3C
      port map(A => \General_Controller_0/uc_rx_byte_0[2]_net_1\, 
        B => \General_Controller_0/uc_rx_byte[7]_net_1\, C => 
        \General_Controller_0/uc_rx_byte[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74116);
    
    HIEFFPLA_INST_0_66877 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73014);
    
    HIEFFPLA_INST_0_58488 : AX1C
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, B => 
        General_Controller_0_en_data_saving, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74752);
    
    \Communications_0/FFU_Command_Checker_0/command_out[0]\ : 
        DFN1E1C1
      port map(D => \Communications_0/UART_0_recv[0]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75625, Q => \Communications_0_ext_recv[0]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[5]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72214, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[5]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[8]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72919, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[8]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_WRITE_RESET_P\ : DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_12_Q\, 
        CLK => CLKINT_0_Y_0, CLR => \AFLSDF_INV_34\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P\);
    
    HIEFFPLA_INST_0_70526 : XOR2
      port map(A => HIEFFPLA_NET_0_72120, B => 
        \Timekeeper_0_milliseconds[7]\, Y => HIEFFPLA_NET_0_72095);
    
    HIEFFPLA_INST_0_61092 : NOR3A
      port map(A => HIEFFPLA_NET_0_74278, B => 
        \Timekeeper_0_milliseconds[17]\, C => 
        \Timekeeper_0_milliseconds[21]\, Y => 
        HIEFFPLA_NET_0_74279);
    
    HIEFFPLA_INST_0_66395 : MX2A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_num_bytes[0]\, 
        S => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_73130);
    
    HIEFFPLA_INST_0_67234 : OR3B
      port map(A => HIEFFPLA_NET_0_72931, B => 
        HIEFFPLA_NET_0_72888, C => HIEFFPLA_NET_0_72883, Y => 
        HIEFFPLA_NET_0_72932);
    
    HIEFFPLA_INST_0_66084 : NOR2A
      port map(A => \Science_0/DAC_SET_0/vector[17]_net_1\, B => 
        \Science_0/DAC_SET_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73214);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[4]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[0]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72777, Q => 
        \Sensors_0_acc_y[4]\);
    
    HIEFFPLA_INST_0_61190 : OR3B
      port map(A => HIEFFPLA_NET_0_74250, B => 
        HIEFFPLA_NET_0_74254, C => HIEFFPLA_NET_0_74244, Y => 
        HIEFFPLA_NET_0_74255);
    
    HIEFFPLA_INST_0_55605 : NAND3
      port map(A => 
        \Communications_0/UART_1/rx_clk_count[29]_net_1\, B => 
        \Communications_0/UART_1/rx_clk_count[30]_net_1\, C => 
        \Communications_0/UART_1/rx_clk_count_c0\, Y => 
        HIEFFPLA_NET_0_75467);
    
    HIEFFPLA_INST_0_68768 : AO1
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[3]_net_1\, C
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72566);
    
    HIEFFPLA_INST_0_66260 : AND2
      port map(A => \Science_0/SET_LP_GAIN_0/state[4]_net_1\, B
         => \Science_0/ADC_READ_0_G4[0]\, Y => 
        HIEFFPLA_NET_0_73163);
    
    HIEFFPLA_INST_0_61103 : NAND3C
      port map(A => \Timekeeper_0_milliseconds[20]\, B => 
        \Timekeeper_0_milliseconds[18]\, C => 
        \Timekeeper_0_milliseconds[12]\, Y => 
        HIEFFPLA_NET_0_74276);
    
    \General_Controller_0/sweep_table_read_value[11]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74168, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[11]_net_1\);
    
    \Communications_0/UART_1/tx_clk_count[2]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75409, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_clk_count_i_0[2]\);
    
    HIEFFPLA_INST_0_70522 : XOR2
      port map(A => HIEFFPLA_NET_0_72117, B => 
        \Timekeeper_0_milliseconds[5]\, Y => HIEFFPLA_NET_0_72097);
    
    HIEFFPLA_INST_0_66129 : NOR2A
      port map(A => \Science_0/DAC_SET_0/vector[12]_net_1\, B => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73200);
    
    HIEFFPLA_INST_0_66380 : AOI1
      port map(A => HIEFFPLA_NET_0_73107, B => 
        HIEFFPLA_NET_0_73038, C => 
        \Sensors_0/Accelerometer_0/state[8]\, Y => 
        HIEFFPLA_NET_0_73134);
    
    \UC_RESET_pad/U0/U0\ : IOPAD_TRI
      port map(D => \UC_RESET_pad/U0/NET1\, E => 
        \UC_RESET_pad/U0/NET2\, PAD => UC_RESET);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[2]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[2]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[2]\);
    
    HIEFFPLA_INST_0_67690 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[6]_net_1\, 
        B => HIEFFPLA_NET_0_72778, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72823);
    
    HIEFFPLA_INST_0_55917 : NOR3B
      port map(A => HIEFFPLA_NET_0_75394, B => 
        \Communications_0/UART_1/tx_count[0]_net_1\, C => 
        HIEFFPLA_NET_0_75420, Y => HIEFFPLA_NET_0_75395);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[17]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72282, Q => 
        \Sensors_0_pressure_temp_raw[17]\);
    
    HIEFFPLA_INST_0_70966 : AO1
      port map(A => HIEFFPLA_NET_0_72000, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        C => HIEFFPLA_NET_0_73150, Y => HIEFFPLA_NET_0_73147);
    
    \Science_0/ADC_READ_0/chan1_data[10]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[10]\);
    
    HIEFFPLA_INST_0_66357 : AX1A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        B => HIEFFPLA_NET_0_73054, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73139);
    
    HIEFFPLA_INST_0_65584 : NOR2A
      port map(A => HIEFFPLA_NET_0_73276, B => 
        \Science_0/ADC_READ_0/cnt3up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73338);
    
    HIEFFPLA_INST_0_61826 : XAI1
      port map(A => Communications_0_uc_rx_rdy, B => 
        \General_Controller_0/uc_rx_state[0]_net_1\, C => 
        HIEFFPLA_NET_0_73943, Y => HIEFFPLA_NET_0_74121);
    
    \Data_Saving_0/Packet_Saver_0/data_out[25]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75219, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[25]\);
    
    HIEFFPLA_INST_0_71129 : AO1
      port map(A => \ch3_data_net_0[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_71977, Y => HIEFFPLA_NET_0_75070);
    
    \Communications_0/UART_0/rx_byte[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75380, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75608, Q => 
        \Communications_0/UART_0/rx_byte[4]_net_1\);
    
    HIEFFPLA_INST_0_66286 : AO1C
      port map(A => HIEFFPLA_NET_0_73171, B => 
        \Science_0/SET_LP_GAIN_0/state[5]_net_1\, C => 
        \Science_0/SET_LP_GAIN_0/state_i_0[1]\, Y => 
        HIEFFPLA_NET_0_73155);
    
    HIEFFPLA_INST_0_71214 : AXOI1
      port map(A => HIEFFPLA_NET_0_75564, B => 
        \Communications_0/UART_0/rx_count[0]_net_1\, C => 
        HIEFFPLA_NET_0_75555, Y => HIEFFPLA_NET_0_71972);
    
    HIEFFPLA_INST_0_56305 : AX1C
      port map(A => HIEFFPLA_NET_0_75308, B => 
        \Data_Saving_0/Packet_Saver_0_we\, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[2]\\\\\, Y
         => HIEFFPLA_NET_0_75312);
    
    \Science_0/ADC_READ_0/cnt2dn[6]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73370, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2dn[6]_net_1\);
    
    HIEFFPLA_INST_0_56332 : AND3A
      port map(A => \Data_Saving_0/FPGA_Buffer_0/full\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[1]\\\\\, C
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[0]\\\\\, 
        Y => HIEFFPLA_NET_0_75308);
    
    \Science_0/ADC_READ_0/cnt[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73282, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73242, Q => 
        \Science_0/ADC_READ_0/cnt[7]_net_1\);
    
    HIEFFPLA_INST_0_56762 : MX2
      port map(A => HIEFFPLA_NET_0_75178, B => 
        HIEFFPLA_NET_0_75035, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75213);
    
    HIEFFPLA_INST_0_56037 : AND2
      port map(A => HIEFFPLA_NET_0_75361, B => 
        HIEFFPLA_NET_0_75326, Y => HIEFFPLA_NET_0_75362);
    
    \ACS_pad/U0/U1\ : IOTRI_OB_EB
      port map(D => ACS_c, E => \VCC\, DOUT => \ACS_pad/U0/NET1\, 
        EOUT => \ACS_pad/U0/NET2\);
    
    \Science_0/ADC_RESET_0/state[0]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73233, CLK => \s_time[5]\, E
         => CLKINT_1_Y, Q => 
        \Science_0/ADC_RESET_0/state[0]_net_1\);
    
    HIEFFPLA_INST_0_68931 : NOR3B
      port map(A => General_Controller_0_en_sensors, B => 
        \Sensors_0/Gyro_0/state[8]\, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, Y
         => HIEFFPLA_NET_0_72518);
    
    HIEFFPLA_INST_0_66754 : NAND2
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\, 
        B => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73045);
    
    HIEFFPLA_INST_0_68166 : AND3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        C => HIEFFPLA_NET_0_72747, Y => HIEFFPLA_NET_0_72718);
    
    HIEFFPLA_INST_0_61261 : AND2A
      port map(A => HIEFFPLA_NET_0_74217, B => 
        HIEFFPLA_NET_0_74233, Y => HIEFFPLA_NET_0_74234);
    
    HIEFFPLA_INST_0_58407 : AO1
      port map(A => \Data_Hub_Packets_0_status_packet[41]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        C => HIEFFPLA_NET_0_75085, Y => HIEFFPLA_NET_0_74776);
    
    \Sensors_0/Gyro_0/I2C_Master_0/data_out[4]\ : DFN0E1C1
      port map(D => GYRO_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72679, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[4]\);
    
    HIEFFPLA_INST_0_57833 : AO1
      port map(A => \Science_0_exp_packet_0[74]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75142, Y => HIEFFPLA_NET_0_74931);
    
    HIEFFPLA_INST_0_56826 : MX2
      port map(A => HIEFFPLA_NET_0_75168, B => 
        HIEFFPLA_NET_0_75019, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75206);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[3]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75264, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\);
    
    HIEFFPLA_INST_0_60883 : NOR3A
      port map(A => \General_Controller_0/command[6]_net_1\, B
         => \General_Controller_0/command[5]_net_1\, C => 
        \General_Controller_0/command[7]_net_1\, Y => 
        HIEFFPLA_NET_0_74331);
    
    HIEFFPLA_INST_0_66057 : AND3
      port map(A => \Science_0/DAC_SET_0/cnt[2]_net_1\, B => 
        \Science_0/DAC_SET_0/cnt[3]_net_1\, C => 
        \Science_0/DAC_SET_0/cnt[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73224);
    
    HIEFFPLA_INST_0_65963 : AOI1B
      port map(A => \Science_0/ADC_READ_0/cnt3up[4]_net_1\, B => 
        HIEFFPLA_NET_0_73276, C => \Science_0/ADC_READ_0_G3[0]\, 
        Y => HIEFFPLA_NET_0_73251);
    
    HIEFFPLA_INST_0_70643 : XA1B
      port map(A => \Timing_0/s_count[1]_net_1\, B => 
        HIEFFPLA_NET_0_72026, C => HIEFFPLA_NET_0_72058, Y => 
        HIEFFPLA_NET_0_72055);
    
    HIEFFPLA_INST_0_64895 : NAND2
      port map(A => HIEFFPLA_NET_0_73514, B => 
        HIEFFPLA_NET_0_73518, Y => HIEFFPLA_NET_0_73515);
    
    HIEFFPLA_INST_0_58017 : AO1B
      port map(A => \Sensors_0_mag_time[17]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74877, Y => HIEFFPLA_NET_0_74878);
    
    HIEFFPLA_INST_0_57269 : AND2
      port map(A => \Sensors_0_mag_time[13]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, Y
         => HIEFFPLA_NET_0_75102);
    
    HIEFFPLA_INST_0_63988 : MX2
      port map(A => HIEFFPLA_NET_0_73653, B => 
        HIEFFPLA_NET_0_73645, S => HIEFFPLA_NET_0_73599, Y => 
        HIEFFPLA_NET_0_73682);
    
    \Data_Saving_0/Packet_Saver_0/data_out[3]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75210, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[3]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[63]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[7]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[63]\);
    
    \General_Controller_0/unit_id[0]\ : DFN1E0P1
      port map(D => \General_Controller_0/uc_rx_byte_0[0]_net_1\, 
        CLK => CLKINT_0_Y_0, PRE => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73990, Q => 
        \General_Controller_0_unit_id[0]\);
    
    \General_Controller_0/uc_rx_prev_state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74059, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_prev_state[0]_net_1\);
    
    HIEFFPLA_INST_0_58298 : AO1
      port map(A => \Sensors_0_acc_x[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74807, Y => HIEFFPLA_NET_0_74808);
    
    HIEFFPLA_INST_0_58103 : AND2
      port map(A => \ch3_data_net_0[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_74854);
    
    HIEFFPLA_INST_0_59943 : MX2
      port map(A => \Science_0_chan1_data[9]\, B => 
        \Science_0_chan0_data[1]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74485);
    
    \Data_Saving_0/Packet_Saver_0/we\ : DFN0E1C1
      port map(D => \Data_Saving_0/Packet_Saver_0/state[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        General_Controller_0_en_data_saving, Q => 
        \Data_Saving_0/Packet_Saver_0_we\);
    
    \Science_0/DAC_SET_0/cnt[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73218, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/cnt[1]_net_1\);
    
    HIEFFPLA_INST_0_56945 : MX2
      port map(A => HIEFFPLA_NET_0_74975, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[8]_net_1\, 
        S => \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, 
        Y => HIEFFPLA_NET_0_75192);
    
    HIEFFPLA_INST_0_67454 : NOR3A
      port map(A => HIEFFPLA_NET_0_72772, B => 
        HIEFFPLA_NET_0_72902, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72875);
    
    HIEFFPLA_INST_0_55533 : NOR2A
      port map(A => \Communications_0/UART_1/rx_count[1]_net_1\, 
        B => \Communications_0/UART_1/rx_count[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75485);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/i2c_addr_1[0]\ : 
        DFN1E0
      port map(D => HIEFFPLA_NET_0_72317, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_72316, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_i2c_addr[0]\);
    
    HIEFFPLA_INST_0_60536 : MX2
      port map(A => \Science_0_chan0_data[6]\, B => 
        \Science_0_chan0_data[10]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74399);
    
    HIEFFPLA_INST_0_70699 : AND2
      port map(A => HIEFFPLA_NET_0_72038, B => \s_time[5]\, Y => 
        HIEFFPLA_NET_0_72039);
    
    HIEFFPLA_INST_0_66708 : AO1
      port map(A => HIEFFPLA_NET_0_73064, B => 
        HIEFFPLA_NET_0_73144, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_73057);
    
    HIEFFPLA_INST_0_67742 : AO1
      port map(A => HIEFFPLA_NET_0_72840, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72811);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[12]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72281, Q => \Sensors_0_pressure_raw[12]\);
    
    HIEFFPLA_INST_0_62821 : AO1
      port map(A => HIEFFPLA_NET_0_73870, B => 
        HIEFFPLA_NET_0_73780, C => HIEFFPLA_NET_0_73992, Y => 
        HIEFFPLA_NET_0_73893);
    
    \General_Controller_0/sweep_table_read_value[9]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74155, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[9]_net_1\);
    
    HIEFFPLA_INST_0_57457 : AO1
      port map(A => \Sensors_0_acc_z[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[12]_net_1\, 
        C => HIEFFPLA_NET_0_74865, Y => HIEFFPLA_NET_0_75040);
    
    HIEFFPLA_INST_0_64609 : NOR3B
      port map(A => \General_Controller_0/uc_tx_state[4]_net_1\, 
        B => \General_Controller_0/uc_tx_substate[1]_net_1\, C
         => HIEFFPLA_NET_0_73563, Y => HIEFFPLA_NET_0_73589);
    
    HIEFFPLA_INST_0_58857 : AND3C
      port map(A => HIEFFPLA_NET_0_74671, B => 
        HIEFFPLA_NET_0_74371, C => HIEFFPLA_NET_0_74552, Y => 
        HIEFFPLA_NET_0_74672);
    
    HIEFFPLA_INST_0_58930 : AND3
      port map(A => HIEFFPLA_NET_0_74568, B => 
        HIEFFPLA_NET_0_74574, C => HIEFFPLA_NET_0_74652, Y => 
        HIEFFPLA_NET_0_74656);
    
    HIEFFPLA_INST_0_59727 : MX2
      port map(A => HIEFFPLA_NET_0_74537, B => 
        HIEFFPLA_NET_0_74523, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74516);
    
    \Data_Saving_0/Packet_Saver_0/data_out[5]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75208, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[5]\);
    
    HIEFFPLA_INST_0_56572 : MX2
      port map(A => HIEFFPLA_NET_0_75203, B => 
        HIEFFPLA_NET_0_75079, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75236);
    
    HIEFFPLA_INST_0_66334 : NAND3
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73143);
    
    \Science_0/ADC_READ_0/exp_packet_1[76]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[20]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[76]\);
    
    HIEFFPLA_INST_0_59917 : MX2
      port map(A => \ch3_data_net_0[3]\, B => \ch3_data_net_0[7]\, 
        S => \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74488);
    
    HIEFFPLA_INST_0_69182 : AO1D
      port map(A => HIEFFPLA_NET_0_72492, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        C => HIEFFPLA_NET_0_72447, Y => HIEFFPLA_NET_0_72453);
    
    HIEFFPLA_INST_0_57169 : AND2
      port map(A => \Sensors_0_pressure_time[18]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75141);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[8]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72281, Q => \Sensors_0_pressure_raw[8]\);
    
    HIEFFPLA_INST_0_57153 : AND2
      port map(A => \Sensors_0_pressure_time[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, Y
         => HIEFFPLA_NET_0_75152);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[22]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[22]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[22]\);
    
    HIEFFPLA_INST_0_65588 : NOR3A
      port map(A => HIEFFPLA_NET_0_73276, B => 
        \Science_0/ADC_READ_0/cnt3up[0]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt3up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73336);
    
    HIEFFPLA_INST_0_67410 : OR3A
      port map(A => HIEFFPLA_NET_0_72911, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[1]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72888);
    
    HIEFFPLA_INST_0_55226 : MX2A
      port map(A => HIEFFPLA_NET_0_75556, B => 
        HIEFFPLA_NET_0_75553, S => 
        \Communications_0/UART_0/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75557);
    
    HIEFFPLA_INST_0_60328 : MX2
      port map(A => HIEFFPLA_NET_0_74473, B => 
        HIEFFPLA_NET_0_74494, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74431);
    
    HIEFFPLA_INST_0_58790 : AO1
      port map(A => HIEFFPLA_NET_0_74405, B => 
        HIEFFPLA_NET_0_74633, C => HIEFFPLA_NET_0_74683, Y => 
        HIEFFPLA_NET_0_74684);
    
    HIEFFPLA_INST_0_58306 : AO1
      port map(A => \Sensors_0_acc_y[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74805, Y => HIEFFPLA_NET_0_74806);
    
    HIEFFPLA_INST_0_55020 : XOR2
      port map(A => \General_Controller_0_unit_id[4]\, B => 
        \Communications_0/UART_0_recv[4]\, Y => 
        HIEFFPLA_NET_0_75614);
    
    \Science_0/ADC_READ_0/exp_packet_1[48]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[14]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[48]\);
    
    HIEFFPLA_INST_0_66541 : OR3A
      port map(A => ACCE_SCL_c, B => HIEFFPLA_NET_0_73095, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[0]_net_1\, 
        Y => HIEFFPLA_NET_0_73096);
    
    HIEFFPLA_INST_0_61987 : XOR2
      port map(A => \General_Controller_0/uc_rx_byte[3]_net_1\, B
         => \General_Controller_0/uc_rx_byte[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74080);
    
    HIEFFPLA_INST_0_65227 : NAND3A
      port map(A => HIEFFPLA_NET_0_73457, B => 
        \Sensors_0_pressure_raw[7]\, C => 
        \Sensors_0_pressure_raw[5]\, Y => HIEFFPLA_NET_0_73440);
    
    HIEFFPLA_INST_0_69292 : NAND3
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[2]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72427);
    
    HIEFFPLA_INST_0_65742 : AND2B
      port map(A => \Science_0/ADC_READ_0/cnt[0]_net_1\, B => 
        HIEFFPLA_NET_0_73241, Y => HIEFFPLA_NET_0_73292);
    
    HIEFFPLA_INST_0_64387 : MX2
      port map(A => HIEFFPLA_NET_0_73711, B => 
        HIEFFPLA_NET_0_73703, S => HIEFFPLA_NET_0_73593, Y => 
        HIEFFPLA_NET_0_73631);
    
    HIEFFPLA_INST_0_58393 : AO1
      port map(A => \Sensors_0_gyro_x[12]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74780, Y => HIEFFPLA_NET_0_74781);
    
    HIEFFPLA_INST_0_57137 : AND2
      port map(A => \Sensors_0_pressure_temp_raw[17]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        Y => HIEFFPLA_NET_0_75160);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[23]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72282, Q => 
        \Sensors_0_pressure_temp_raw[23]\);
    
    \General_Controller_0/constant_bias_probe_id[7]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73923, Q => 
        \General_Controller_0/un10_uc_tx_rdy_i[7]\);
    
    \Timekeeper_0/old_1kHz\ : DFN1E0
      port map(D => \m_time[7]\, CLK => CLKINT_0_Y_0, E => 
        CLKINT_1_Y, Q => \Timekeeper_0/old_1kHz_net_1\);
    
    HIEFFPLA_INST_0_61921 : NOR3B
      port map(A => HIEFFPLA_NET_0_74076, B => 
        HIEFFPLA_NET_0_74085, C => 
        \General_Controller_0/uc_rx_byte[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74098);
    
    \General_Controller_0/uc_tx_state[3]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73570, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[3]_net_1\);
    
    HIEFFPLA_INST_0_71033 : AO1A
      port map(A => HIEFFPLA_NET_0_73559, B => 
        HIEFFPLA_NET_0_71986, C => HIEFFPLA_NET_0_73590, Y => 
        HIEFFPLA_NET_0_73606);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_y[7]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72783, Q => 
        \Sensors_0_mag_y[7]\);
    
    \Science_0/ADC_READ_0/chan3_data[6]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[12]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[6]\);
    
    HIEFFPLA_INST_0_58258 : AO1
      port map(A => \Sensors_0_gyro_time[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75110, Y => HIEFFPLA_NET_0_74818);
    
    \Communications_0/UART_0/rx_byte[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75380, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75607, Q => 
        \Communications_0/UART_0/rx_byte[5]_net_1\);
    
    HIEFFPLA_INST_0_63297 : XO1A
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, C => 
        HIEFFPLA_NET_0_73786, Y => HIEFFPLA_NET_0_73784);
    
    HIEFFPLA_INST_0_69261 : NAND3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, B
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, 
        C => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, Y => 
        HIEFFPLA_NET_0_72436);
    
    HIEFFPLA_INST_0_63321 : NOR3A
      port map(A => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, B => 
        HIEFFPLA_NET_0_73786, C => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73777);
    
    HIEFFPLA_INST_0_61021 : OA1A
      port map(A => \General_Controller_0/flight_state[1]_net_1\, 
        B => HIEFFPLA_NET_0_74257, C => HIEFFPLA_NET_0_74298, Y
         => HIEFFPLA_NET_0_74293);
    
    HIEFFPLA_INST_0_58772 : NAND3C
      port map(A => HIEFFPLA_NET_0_74674, B => 
        HIEFFPLA_NET_0_74677, C => HIEFFPLA_NET_0_74688, Y => 
        HIEFFPLA_NET_0_74689);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/data_out_1[4]\ : 
        DFN1E0C1
      port map(D => \AFLSDF_INV_35\, CLK => CLKINT_0_Y_0, CLR => 
        CLKINT_1_Y, E => HIEFFPLA_NET_0_72270, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[4]\);
    
    HIEFFPLA_INST_0_61436 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[47]\, B => 
        \Timekeeper_0_milliseconds[7]\, S => HIEFFPLA_NET_0_74266, 
        Y => HIEFFPLA_NET_0_74199);
    
    HIEFFPLA_INST_0_68794 : NAND2B
      port map(A => HIEFFPLA_NET_0_72485, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/isSetup_net_1\, Y
         => HIEFFPLA_NET_0_72559);
    
    HIEFFPLA_INST_0_59689 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[58]\, B => 
        \Data_Hub_Packets_0_status_packet[62]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74522);
    
    HIEFFPLA_INST_0_57759 : AO1B
      port map(A => \Sensors_0_acc_time[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74950, Y => HIEFFPLA_NET_0_74951);
    
    HIEFFPLA_INST_0_67930 : OR3A
      port map(A => HIEFFPLA_NET_0_72919, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        Y => HIEFFPLA_NET_0_72770);
    
    \Data_Saving_0/Packet_Saver_0/data_out[1]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75225, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[1]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[56]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[0]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[56]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[7]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72919, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[7]_net_1\);
    
    HIEFFPLA_INST_0_60839 : NOR3B
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/state[6]_net_1\, C => 
        Communications_0_ext_tx_rdy, Y => HIEFFPLA_NET_0_74348);
    
    \Communications_0/UART_1/rx_clk_count[30]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75457, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75443, Q => 
        \Communications_0/UART_1/rx_clk_count[30]_net_1\);
    
    HIEFFPLA_INST_0_57867 : AO1B
      port map(A => \Sensors_0_mag_time[22]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_74920, Y => HIEFFPLA_NET_0_74921);
    
    \Science_0/ADC_READ_0/cnt3dn[5]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73342, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73423, Q => 
        \Science_0/ADC_READ_0/cnt3dn[5]_net_1\);
    
    HIEFFPLA_INST_0_55698 : AND2
      port map(A => \Communications_0/UART_1/rx_state[0]_net_1\, 
        B => \Communications_0/UART_1/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75444);
    
    \Science_0/ADC_READ_0/exp_packet_1[40]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[6]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[40]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[5]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72279, Q => 
        \Sensors_0_pressure_temp_raw[5]\);
    
    HIEFFPLA_INST_0_62539 : OA1C
      port map(A => HIEFFPLA_NET_0_73856, B => 
        HIEFFPLA_NET_0_73811, C => HIEFFPLA_NET_0_73955, Y => 
        HIEFFPLA_NET_0_73961);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_4\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[4]\\\\\, CLK => 
        CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_4_Q\);
    
    HIEFFPLA_INST_0_70381 : AND3
      port map(A => \Timekeeper_0_microseconds[11]\, B => 
        HIEFFPLA_NET_0_72152, C => 
        \Timekeeper_0_microseconds[12]\, Y => 
        HIEFFPLA_NET_0_72155);
    
    HIEFFPLA_INST_0_65725 : NAND2B
      port map(A => \Science_0/ADC_READ_0/cnt[5]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73298);
    
    HIEFFPLA_INST_0_55885 : AX1B
      port map(A => \Communications_0/UART_1/tx_clk_count_i_0[5]\, 
        B => HIEFFPLA_NET_0_75412, C => 
        \Communications_0/UART_1/tx_clk_count_i_0[6]\, Y => 
        HIEFFPLA_NET_0_75404);
    
    HIEFFPLA_INST_0_55155 : XA1B
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[26]_net_1\, B => 
        HIEFFPLA_NET_0_75586, C => HIEFFPLA_NET_0_75567, Y => 
        HIEFFPLA_NET_0_75573);
    
    HIEFFPLA_INST_0_65978 : OA1C
      port map(A => HIEFFPLA_NET_0_73246, B => 
        \Science_0/ADC_READ_0_G4[1]\, C => HIEFFPLA_NET_0_73319, 
        Y => HIEFFPLA_NET_0_73248);
    
    \Science_0/ADC_READ_0/data_a[12]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_a[12]_net_1\);
    
    \General_Controller_0/state_seconds[7]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74220, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[7]_net_1\);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72416, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[3]_net_1\);
    
    HIEFFPLA_INST_0_69657 : MX2
      port map(A => HIEFFPLA_NET_0_72425, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        S => PRESSURE_SCL_c, Y => HIEFFPLA_NET_0_72335);
    
    HIEFFPLA_INST_0_65858 : MX2
      port map(A => \Science_0/ADC_READ_0_G1[1]\, B => 
        \Science_0/ADC_READ_0_G3[1]\, S => 
        \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73269);
    
    HIEFFPLA_INST_0_58389 : AO1
      port map(A => \Sensors_0_mag_x[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_75107, Y => HIEFFPLA_NET_0_74782);
    
    \Communications_0/UART_0/recv[7]\ : DFN1E1C1
      port map(D => \Communications_0/UART_0/rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75551, Q => 
        \Communications_0/UART_0_recv[7]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[6]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72503, Q => 
        \Sensors_0_gyro_x[6]\);
    
    \General_Controller_0/st_wdata[4]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[4]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[9]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72283, Q => 
        \Sensors_0_pressure_temp_raw[9]\);
    
    HIEFFPLA_INST_0_61606 : AND3
      port map(A => HIEFFPLA_NET_0_73778, B => 
        HIEFFPLA_NET_0_74173, C => HIEFFPLA_NET_0_73972, Y => 
        HIEFFPLA_NET_0_74175);
    
    \Science_0/ADC_READ_0/chan4_data[5]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan4_data[5]\);
    
    HIEFFPLA_INST_0_58750 : AND3
      port map(A => \GS_Readout_0/state[3]_net_1\, B => 
        HIEFFPLA_NET_0_74372, C => HIEFFPLA_NET_0_74552, Y => 
        HIEFFPLA_NET_0_74693);
    
    HIEFFPLA_INST_0_61087 : NOR3A
      port map(A => HIEFFPLA_NET_0_74279, B => 
        HIEFFPLA_NET_0_74276, C => 
        \Timekeeper_0_milliseconds[22]\, Y => 
        HIEFFPLA_NET_0_74280);
    
    HIEFFPLA_INST_0_56397 : NOR3B
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, B
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, 
        C => HIEFFPLA_NET_0_75370, Y => HIEFFPLA_NET_0_75290);
    
    HIEFFPLA_INST_0_59897 : MX2
      port map(A => HIEFFPLA_NET_0_74395, B => 
        HIEFFPLA_NET_0_74407, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74490);
    
    \Timekeeper_0/microseconds[18]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72142, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[18]\);
    
    AFLSDF_INV_11 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_11\);
    
    HIEFFPLA_INST_0_64585 : NOR2A
      port map(A => HIEFFPLA_NET_0_73602, B => 
        HIEFFPLA_NET_0_73938, Y => HIEFFPLA_NET_0_73595);
    
    HIEFFPLA_INST_0_60302 : MX2
      port map(A => \Science_0_chan5_data[2]\, B => 
        \Science_0_chan5_data[6]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74434);
    
    HIEFFPLA_INST_0_69857 : NAND2B
      port map(A => \Sensors_0/Pressure_Sensor_0/state[8]\, B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_num_bytes[0]\, 
        Y => HIEFFPLA_NET_0_72289);
    
    HIEFFPLA_INST_0_56745 : AOI1B
      port map(A => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[1]_net_1\, B => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, C => 
        HIEFFPLA_NET_0_75183, Y => HIEFFPLA_NET_0_75217);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72866, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72864, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\);
    
    HIEFFPLA_INST_0_60610 : AND2B
      port map(A => \GS_Readout_0/subState[0]_net_1\, B => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74387);
    
    HIEFFPLA_INST_0_60485 : AND3
      port map(A => HIEFFPLA_NET_0_74341, B => 
        HIEFFPLA_NET_0_74342, C => HIEFFPLA_NET_0_74560, Y => 
        HIEFFPLA_NET_0_74407);
    
    \Communications_0/UART_0/rx_clk_count[26]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75573, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75554, Q => 
        \Communications_0/UART_0/rx_clk_count[26]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72468, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[1]_net_1\);
    
    \GS_Readout_0/state[5]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74601, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \GS_Readout_0/state[5]_net_1\);
    
    \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/we\ : 
        DFN1E0C1
      port map(D => HIEFFPLA_NET_0_72173, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72172, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_we\);
    
    HIEFFPLA_INST_0_66268 : NAND2
      port map(A => HIEFFPLA_NET_0_73166, B => 
        \Science_0/SET_LP_GAIN_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73161);
    
    HIEFFPLA_INST_0_61972 : AND3
      port map(A => HIEFFPLA_NET_0_74106, B => 
        HIEFFPLA_NET_0_74077, C => HIEFFPLA_NET_0_74073, Y => 
        HIEFFPLA_NET_0_74086);
    
    \Communications_0/UART_0/tx_rdy\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75501, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => Communications_0_ext_tx_rdy);
    
    HIEFFPLA_INST_0_68883 : NAND3B
      port map(A => HIEFFPLA_NET_0_72513, B => 
        HIEFFPLA_NET_0_72517, C => HIEFFPLA_NET_0_72532, Y => 
        HIEFFPLA_NET_0_72533);
    
    HIEFFPLA_INST_0_64437 : MX2
      port map(A => HIEFFPLA_NET_0_73706, B => 
        HIEFFPLA_NET_0_73698, S => HIEFFPLA_NET_0_73593, Y => 
        HIEFFPLA_NET_0_73626);
    
    HIEFFPLA_INST_0_63014 : NAND3C
      port map(A => \General_Controller_0/uc_rx_byte[0]_net_1\, B
         => HIEFFPLA_NET_0_74082, C => 
        \General_Controller_0/uc_rx_byte[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73847);
    
    \ClockDivs_0/clk_800kHz_RNIT3EB\ : CLKINT
      port map(A => \ClockDivs_0/clk_800kHz_i\, Y => 
        ClockDivs_0_clk_800kHz);
    
    HIEFFPLA_INST_0_71009 : NAND3
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[2]_net_1\, 
        B => \Pressure_Signal_Debounce_0/ms_cnt[3]_net_1\, C => 
        \Pressure_Signal_Debounce_0/ms_cnt[1]_net_1\, Y => 
        HIEFFPLA_NET_0_71991);
    
    \General_Controller_0/constant_bias_voltage_1[2]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[2]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74321, Q => 
        \General_Controller_0/constant_bias_voltage_1[2]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/data_out[0]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75236, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[0]\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/data_out[7]\ : DFN0E1C1
      port map(D => GYRO_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72673, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[7]\);
    
    \Science_0/ADC_READ_0/cnt4up[4]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73301, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4up[4]_net_1\);
    
    HIEFFPLA_INST_0_70428 : XOR2
      port map(A => HIEFFPLA_NET_0_72154, B => 
        \Timekeeper_0_microseconds[3]\, Y => HIEFFPLA_NET_0_72134);
    
    HIEFFPLA_INST_0_61026 : AO1A
      port map(A => HIEFFPLA_NET_0_74257, B => 
        \General_Controller_0/flight_state[1]_net_1\, C => 
        \General_Controller_0/flight_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74292);
    
    HIEFFPLA_INST_0_65864 : MX2
      port map(A => \Science_0/ADC_READ_0_G2[0]\, B => 
        \Science_0/ADC_READ_0_G4[0]\, S => 
        \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73268);
    
    HIEFFPLA_INST_0_67967 : NAND3C
      port map(A => HIEFFPLA_NET_0_72738, B => 
        HIEFFPLA_NET_0_72717, C => HIEFFPLA_NET_0_72744, Y => 
        HIEFFPLA_NET_0_72765);
    
    \Communications_0/UART_0/tx_byte[2]\ : DFN1E1
      port map(D => \GS_Readout_0_send[2]\, CLK => CLKINT_0_Y_0, 
        E => HIEFFPLA_NET_0_75504, Q => 
        \Communications_0/UART_0/tx_byte[2]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[12]\ : DFN1E0
      port map(D => \AFLSDF_INV_36\, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_73243, Q => \Science_0_exp_packet_0[12]\);
    
    HIEFFPLA_INST_0_63310 : AND2
      port map(A => 
        \General_Controller_0/uc_rx_substate[0]_net_1\, B => 
        \General_Controller_0/uc_rx_substate[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73780);
    
    HIEFFPLA_INST_0_62262 : AND2B
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74018);
    
    \General_Controller_0/st_wdata[1]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[1]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[1]\);
    
    HIEFFPLA_INST_0_62209 : AXO2
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[3]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74029);
    
    HIEFFPLA_INST_0_70997 : AO1B
      port map(A => \Science_0/ADC_READ_0/cnt1up[4]_net_1\, B => 
        HIEFFPLA_NET_0_73276, C => \Science_0/ADC_READ_0_G1[0]\, 
        Y => HIEFFPLA_NET_0_71994);
    
    HIEFFPLA_INST_0_60848 : AND2
      port map(A => \GS_Readout_0/subState[1]_net_1\, B => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74344);
    
    HIEFFPLA_INST_0_67861 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, B
         => HIEFFPLA_NET_0_72747, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72785);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_time[12]\ : DFN1E1
      port map(D => \Timekeeper_0_microseconds[12]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72546, Q => 
        \Sensors_0_gyro_time[12]\);
    
    HIEFFPLA_INST_0_63566 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[13]_net_1\, B
         => \General_Controller_0/sweep_table_points[13]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73748);
    
    HIEFFPLA_INST_0_61142 : NOR2A
      port map(A => HIEFFPLA_NET_0_74326, B => 
        HIEFFPLA_NET_0_74330, Y => HIEFFPLA_NET_0_74265);
    
    HIEFFPLA_INST_0_55702 : XA1B
      port map(A => \Communications_0/UART_1/rx_state[0]_net_1\, 
        B => \Communications_0/UART_1/rx_state[1]_net_1\, C => 
        HIEFFPLA_NET_0_75482, Y => HIEFFPLA_NET_0_75442);
    
    HIEFFPLA_INST_0_65053 : AOI1D
      port map(A => HIEFFPLA_NET_0_73454, B => 
        HIEFFPLA_NET_0_73453, C => 
        \Pressure_Signal_Debounce_0/state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73480);
    
    HIEFFPLA_INST_0_55265 : MX2
      port map(A => HIEFFPLA_NET_0_75547, B => 
        HIEFFPLA_NET_0_75546, S => 
        \Communications_0/UART_0/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75549);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/temp[0]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[0]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72555, Q => 
        \Sensors_0_gyro_temp[0]\);
    
    HIEFFPLA_INST_0_65715 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt4up[4]_net_1\, B => 
        HIEFFPLA_NET_0_73300, C => HIEFFPLA_NET_0_73309, Y => 
        HIEFFPLA_NET_0_73301);
    
    HIEFFPLA_INST_0_67524 : AO1A
      port map(A => HIEFFPLA_NET_0_72832, B => 
        HIEFFPLA_NET_0_72743, C => HIEFFPLA_NET_0_72823, Y => 
        HIEFFPLA_NET_0_72858);
    
    \General_Controller_0/uc_rx_state_0[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73997, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_rx_state_0[1]_net_1\);
    
    \General_Controller_0/state_seconds[15]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74234, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[15]_net_1\);
    
    \Communications_0/UART_0/tx_byte[0]\ : DFN1E1
      port map(D => \GS_Readout_0_send[0]\, CLK => CLKINT_0_Y_0, 
        E => HIEFFPLA_NET_0_75504, Q => 
        \Communications_0/UART_0/tx_byte[0]_net_1\);
    
    HIEFFPLA_INST_0_62845 : NAND3
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        \General_Controller_0/uc_rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73884);
    
    HIEFFPLA_INST_0_58108 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_74852);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[1]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72804, Q => 
        \Sensors_0_mag_x[1]\);
    
    \Data_Saving_0/Packet_Saver_0/packet_select_1[11]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74772, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\);
    
    \Timekeeper_0/microseconds[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72133, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[4]\);
    
    HIEFFPLA_INST_0_62513 : AO1
      port map(A => HIEFFPLA_NET_0_73805, B => 
        HIEFFPLA_NET_0_73860, C => HIEFFPLA_NET_0_73966, Y => 
        HIEFFPLA_NET_0_73967);
    
    \FMC_DA_pad[2]/U0/U0\ : IOPAD_TRI
      port map(D => \FMC_DA_pad[2]/U0/NET1\, E => 
        \FMC_DA_pad[2]/U0/NET2\, PAD => FMC_DA(2));
    
    \Science_0/ADC_READ_0/exp_packet_1[74]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[18]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[74]\);
    
    HIEFFPLA_INST_0_64998 : AO1B
      port map(A => HIEFFPLA_NET_0_73451, B => 
        HIEFFPLA_NET_0_73477, C => HIEFFPLA_NET_0_73482, Y => 
        HIEFFPLA_NET_0_73492);
    
    HIEFFPLA_INST_0_57499 : AO1B
      port map(A => \Sensors_0_mag_z[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[11]_net_1\, 
        C => HIEFFPLA_NET_0_75027, Y => HIEFFPLA_NET_0_75028);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/data_out[7]\ : 
        DFN0E1C1
      port map(D => ACCE_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73115, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\);
    
    HIEFFPLA_INST_0_66557 : NAND3C
      port map(A => HIEFFPLA_NET_0_73081, B => 
        HIEFFPLA_NET_0_73079, C => 
        \Sensors_0/Accelerometer_0/state_0[8]\, Y => 
        HIEFFPLA_NET_0_73092);
    
    HIEFFPLA_INST_0_59216 : OA1A
      port map(A => HIEFFPLA_NET_0_74382, B => 
        \GS_Readout_0/state[2]_net_1\, C => HIEFFPLA_NET_0_74581, 
        Y => HIEFFPLA_NET_0_74586);
    
    HIEFFPLA_INST_0_57164 : AO1
      port map(A => \Sensors_0_acc_x[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y
         => HIEFFPLA_NET_0_75143);
    
    \Communications_0/UART_1/tx_count[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75393, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75388, Q => 
        \Communications_0/UART_1/tx_count[0]_net_1\);
    
    HIEFFPLA_INST_0_68678 : NAND3C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[3]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_72591);
    
    HIEFFPLA_INST_0_69891 : AND2B
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72277);
    
    HIEFFPLA_INST_0_62711 : NOR3A
      port map(A => HIEFFPLA_NET_0_73860, B => 
        HIEFFPLA_NET_0_73916, C => HIEFFPLA_NET_0_73776, Y => 
        HIEFFPLA_NET_0_73923);
    
    HIEFFPLA_INST_0_70790 : OA1A
      port map(A => HIEFFPLA_NET_0_72012, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/bitcnt[1]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[5]_net_1\, 
        Y => HIEFFPLA_NET_0_72377);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_1\ : DFN0E0P1
      port map(D => HIEFFPLA_NET_0_73073, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73100, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/sda_cl_1_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_y[11]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[7]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72777, Q => 
        \Sensors_0_acc_y[11]\);
    
    HIEFFPLA_INST_0_68812 : NAND2B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[0]_net_1\, B
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0/state[1]_net_1\, 
        Y => HIEFFPLA_NET_0_72551);
    
    HIEFFPLA_INST_0_57671 : AO1
      port map(A => \Sensors_0_pressure_raw[17]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, C
         => HIEFFPLA_NET_0_74974, Y => HIEFFPLA_NET_0_74975);
    
    HIEFFPLA_INST_0_57552 : AOI1
      port map(A => \Science_0_exp_packet_0[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[5]_net_1\, 
        C => HIEFFPLA_NET_0_75011, Y => HIEFFPLA_NET_0_75012);
    
    \Science_0/ADC_READ_0/cnt2up[3]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73361, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2up[3]_net_1\);
    
    HIEFFPLA_INST_0_65373 : NOR3A
      port map(A => HIEFFPLA_NET_0_73276, B => 
        \Science_0/ADC_READ_0/cnt1up[0]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt1up[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73397);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_z[6]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72753, Q => 
        \Sensors_0_acc_z[6]\);
    
    HIEFFPLA_INST_0_69262 : NOR2A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        B => \Sensors_0/Gyro_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72435);
    
    HIEFFPLA_INST_0_67764 : NOR3A
      port map(A => HIEFFPLA_NET_0_72738, B => 
        HIEFFPLA_NET_0_72874, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72807);
    
    HIEFFPLA_INST_0_57158 : AND2
      port map(A => \Sensors_0_pressure_time[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[10]_net_1\, Y
         => HIEFFPLA_NET_0_75147);
    
    HIEFFPLA_INST_0_64951 : XOR2
      port map(A => \I2C_PassThrough_0/cnt[0]_net_1\, B => 
        HIEFFPLA_NET_0_73514, Y => HIEFFPLA_NET_0_73505);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[19]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[19]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[19]\);
    
    HIEFFPLA_INST_0_59194 : NOR2A
      port map(A => \GS_Readout_0/state[5]_net_1\, B => 
        HIEFFPLA_NET_0_74374, Y => HIEFFPLA_NET_0_74591);
    
    HIEFFPLA_INST_0_58944 : NOR2A
      port map(A => \GS_Readout_0/state[2]_net_1\, B => 
        HIEFFPLA_NET_0_74421, Y => HIEFFPLA_NET_0_74652);
    
    \Science_0/ADC_READ_0/data_b[0]\ : DFN1E1C1
      port map(D => AA_c, CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, 
        E => \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[0]_net_1\);
    
    HIEFFPLA_INST_0_61651 : MX2
      port map(A => \SweepTable_0_RD[13]\, B => 
        \SweepTable_1_RD[13]\, S => 
        \General_Controller_0/sweep_table_probe_id[0]_net_1\, Y
         => HIEFFPLA_NET_0_74166);
    
    \Data_Saving_0/Packet_Saver_0/data_out[11]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75234, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[11]\);
    
    \Communications_0/UART_0/tx_clk_count[5]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75521, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_0/tx_clk_count_i_0[5]\);
    
    \Sensors_0/Gyro_0/I2C_Master_0/state[7]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72607, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\);
    
    \Science_0/SET_LP_GAIN_0/state[5]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73154, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/state[5]_net_1\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[2]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[2]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72919, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[2]_net_1\);
    
    HIEFFPLA_INST_0_69902 : NAND2B
      port map(A => HIEFFPLA_NET_0_72269, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out_rdy\, 
        Y => HIEFFPLA_NET_0_72271);
    
    HIEFFPLA_INST_0_55079 : AND3C
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[25]_net_1\, B => 
        \Communications_0/UART_0/rx_clk_count[26]_net_1\, C => 
        \Communications_0/UART_0/rx_clk_count[27]_net_1\, Y => 
        HIEFFPLA_NET_0_75596);
    
    HIEFFPLA_INST_0_70340 : AOI1D
      port map(A => General_Controller_0_st_ren1, B => 
        \SweepTable_0/WEBP\, C => 
        \General_Controller_0_st_raddr_1[2]\, Y => 
        \TableSelect_0_RADDR[2]\);
    
    HIEFFPLA_INST_0_63872 : MX2
      port map(A => HIEFFPLA_NET_0_73670, B => 
        HIEFFPLA_NET_0_73665, S => HIEFFPLA_NET_0_73594, Y => 
        HIEFFPLA_NET_0_73697);
    
    HIEFFPLA_INST_0_64051 : MX2
      port map(A => HIEFFPLA_NET_0_73639, B => 
        HIEFFPLA_NET_0_73631, S => HIEFFPLA_NET_0_73585, Y => 
        HIEFFPLA_NET_0_73676);
    
    HIEFFPLA_INST_0_62682 : NAND3C
      port map(A => HIEFFPLA_NET_0_74028, B => 
        HIEFFPLA_NET_0_73947, C => HIEFFPLA_NET_0_73865, Y => 
        HIEFFPLA_NET_0_73929);
    
    \General_Controller_0/sweep_table_sweep_cnt[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74136, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73927, Q => 
        \General_Controller_0/sweep_table_sweep_cnt[2]_net_1\);
    
    HIEFFPLA_INST_0_68540 : AND3C
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_72622);
    
    HIEFFPLA_INST_0_62071 : AO1A
      port map(A => HIEFFPLA_NET_0_73862, B => 
        HIEFFPLA_NET_0_73916, C => HIEFFPLA_NET_0_74050, Y => 
        HIEFFPLA_NET_0_74058);
    
    HIEFFPLA_INST_0_61796 : NAND2
      port map(A => HIEFFPLA_NET_0_74147, B => 
        \General_Controller_0/sweep_table_sweep_cnt[14]_net_1\, Y
         => HIEFFPLA_NET_0_74128);
    
    HIEFFPLA_INST_0_58890 : AND2
      port map(A => \General_Controller_0_gs_id[0]\, B => 
        HIEFFPLA_NET_0_74484, Y => HIEFFPLA_NET_0_74664);
    
    \General_Controller_0/uc_tx_nextstate[2]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73915, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73857, Q => 
        \General_Controller_0/uc_tx_nextstate[2]_net_1\);
    
    \Science_0/ADC_READ_0/CS\ : DFN1E1P1
      port map(D => \Science_0/ADC_READ_0/countere\, CLK => 
        CLKINT_0_Y_0, PRE => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73425, Q => ACS_c);
    
    HIEFFPLA_INST_0_62657 : NAND3C
      port map(A => HIEFFPLA_NET_0_73897, B => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, C => 
        \General_Controller_0/uc_rx_state_0[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73934);
    
    HIEFFPLA_INST_0_60975 : AND2
      port map(A => \Timekeeper_0_milliseconds[2]\, B => 
        \General_Controller_0/flight_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74306);
    
    \Timing_0/s_time[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72048, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_time[0]_net_1\);
    
    HIEFFPLA_INST_0_62655 : OR3B
      port map(A => HIEFFPLA_NET_0_74010, B => 
        \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73935);
    
    HIEFFPLA_INST_0_67215 : AO1A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_s_ack_error\, B
         => HIEFFPLA_NET_0_72880, C => HIEFFPLA_NET_0_72936, Y
         => HIEFFPLA_NET_0_72937);
    
    HIEFFPLA_INST_0_60639 : OR3A
      port map(A => \GS_Readout_0/subState[4]_net_1\, B => 
        HIEFFPLA_NET_0_74374, C => 
        \GS_Readout_0/subState[1]_net_1\, Y => 
        HIEFFPLA_NET_0_74382);
    
    HIEFFPLA_INST_0_59781 : MX2
      port map(A => \Sensors_0_acc_z[4]\, B => 
        \Sensors_0_acc_z[8]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74509);
    
    \Data_Saving_0/Packet_Saver_0/mag_flag\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_74770, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => 
        General_Controller_0_en_data_saving, Q => 
        \Data_Saving_0/Packet_Saver_0/mag_flag_net_1\);
    
    HIEFFPLA_INST_0_70176 : NOR3B
      port map(A => \Sensors_0/Pressure_Sensor_0/state[8]\, B => 
        HIEFFPLA_NET_0_72278, C => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        Y => HIEFFPLA_NET_0_72201);
    
    HIEFFPLA_INST_0_62442 : NOR3B
      port map(A => HIEFFPLA_NET_0_73900, B => 
        HIEFFPLA_NET_0_73800, C => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73981);
    
    HIEFFPLA_INST_0_62289 : OA1C
      port map(A => HIEFFPLA_NET_0_74025, B => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, C => 
        HIEFFPLA_NET_0_74041, Y => HIEFFPLA_NET_0_74014);
    
    HIEFFPLA_INST_0_60069 : MX2
      port map(A => \ch3_data_net_0[10]\, B => 
        \Sensors_0_acc_z[2]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74466);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[4]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72804, Q => 
        \Sensors_0_mag_x[4]\);
    
    \Science_0/ADC_READ_0/exp_packet_1[54]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/chan[0]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[54]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[4]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[4]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72919, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[4]_net_1\);
    
    HIEFFPLA_INST_0_66919 : NAND3B
      port map(A => HIEFFPLA_NET_0_72929, B => 
        HIEFFPLA_NET_0_72789, C => HIEFFPLA_NET_0_72998, Y => 
        HIEFFPLA_NET_0_73005);
    
    HIEFFPLA_INST_0_67828 : OR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out_rdy\, B
         => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72792);
    
    \Science_0/SET_LP_GAIN_0/state[1]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_73156, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Science_0/SET_LP_GAIN_0/state_i_0[1]\);
    
    \General_Controller_0/st_waddr[2]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_step_id[2]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_waddr[2]\);
    
    \Science_0/ADC_READ_0/cnt1up[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73394, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73418, Q => 
        \Science_0/ADC_READ_0/cnt1up[2]_net_1\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_y[5]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72482, Q => 
        \Sensors_0_gyro_y[5]\);
    
    HIEFFPLA_INST_0_65335 : XA1B
      port map(A => HIEFFPLA_NET_0_73409, B => 
        \Science_0/ADC_READ_0/cnt1dn[2]_net_1\, C => 
        HIEFFPLA_NET_0_73244, Y => HIEFFPLA_NET_0_73406);
    
    HIEFFPLA_INST_0_61967 : AO1A
      port map(A => HIEFFPLA_NET_0_74112, B => 
        HIEFFPLA_NET_0_74074, C => HIEFFPLA_NET_0_74086, Y => 
        HIEFFPLA_NET_0_74087);
    
    HIEFFPLA_INST_0_70723 : AND3
      port map(A => HIEFFPLA_NET_0_72032, B => 
        \Timing_0/m_count[3]_net_1\, C => 
        \Timing_0/m_count[4]_net_1\, Y => HIEFFPLA_NET_0_72031);
    
    \Communications_0/UART_1/recv[6]\ : DFN1E1C1
      port map(D => \Communications_0/UART_1/rx_byte[6]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75441, Q => \Communications_0_uc_recv[6]\);
    
    HIEFFPLA_INST_0_55991 : XA1A
      port map(A => HIEFFPLA_NET_0_75320, B => 
        HIEFFPLA_NET_0_75304, C => HIEFFPLA_NET_0_75374, Y => 
        HIEFFPLA_NET_0_75375);
    
    HIEFFPLA_INST_0_59633 : MX2
      port map(A => HIEFFPLA_NET_0_74536, B => 
        HIEFFPLA_NET_0_74534, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74528);
    
    HIEFFPLA_INST_0_55901 : AXOI4
      port map(A => HIEFFPLA_NET_0_75386, B => 
        \Communications_0/UART_1/tx_clk_count[0]_net_1\, C => 
        \Communications_0/UART_1/tx_clk_count[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75401);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]\ : 
        DFN1P1
      port map(D => HIEFFPLA_NET_0_72856, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[8]_net_1\);
    
    HIEFFPLA_INST_0_67330 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        C => \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        Y => HIEFFPLA_NET_0_72906);
    
    HIEFFPLA_INST_0_55180 : OA1C
      port map(A => \Communications_0/UART_0/rx_state[1]_net_1\, 
        B => HIEFFPLA_NET_0_75552, C => HIEFFPLA_NET_0_75594, Y
         => HIEFFPLA_NET_0_75567);
    
    HIEFFPLA_INST_0_62527 : NOR2A
      port map(A => HIEFFPLA_NET_0_74113, B => 
        HIEFFPLA_NET_0_73963, Y => HIEFFPLA_NET_0_73964);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/num_bytes_1[1]\ : 
        DFN1E0C1
      port map(D => HIEFFPLA_NET_0_72290, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72232, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_num_bytes[1]\);
    
    HIEFFPLA_INST_0_67487 : AO1A
      port map(A => HIEFFPLA_NET_0_72941, B => 
        HIEFFPLA_NET_0_72957, C => HIEFFPLA_NET_0_72835, Y => 
        HIEFFPLA_NET_0_72867);
    
    HIEFFPLA_INST_0_70454 : AND3
      port map(A => \Timekeeper_0_milliseconds[7]\, B => 
        HIEFFPLA_NET_0_72120, C => \Timekeeper_0_milliseconds[8]\, 
        Y => HIEFFPLA_NET_0_72124);
    
    HIEFFPLA_INST_0_58935 : NAND2B
      port map(A => HIEFFPLA_NET_0_74651, B => 
        HIEFFPLA_NET_0_74621, Y => HIEFFPLA_NET_0_74655);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72470, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[11]_net_1\);
    
    HIEFFPLA_INST_0_70807 : AND3B
      port map(A => HIEFFPLA_NET_0_72008, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]_net_1\, 
        C => HIEFFPLA_NET_0_72495, Y => HIEFFPLA_NET_0_72500);
    
    \FMC_CLK_pad/U0/U0\ : IOPAD_IN
      port map(PAD => FMC_CLK, Y => \FMC_CLK_pad/U0/NET1\);
    
    HIEFFPLA_INST_0_60171 : MX2
      port map(A => HIEFFPLA_NET_0_74379, B => 
        HIEFFPLA_NET_0_74377, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74450);
    
    HIEFFPLA_INST_0_59535 : MX2
      port map(A => HIEFFPLA_NET_0_74411, B => 
        HIEFFPLA_NET_0_74430, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74541);
    
    \General_Controller_0/state_seconds[8]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_74219, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74268, Q => 
        \General_Controller_0/state_seconds[8]_net_1\);
    
    \Communications_0/UART_1/tx_byte[3]\ : DFN1E1
      port map(D => \General_Controller_0_uc_send[3]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_75385, Q => 
        \Communications_0/UART_1/tx_byte[3]_net_1\);
    
    HIEFFPLA_INST_0_55487 : AX1
      port map(A => HIEFFPLA_NET_0_75528, B => 
        \Communications_0/UART_0/tx_state[0]_net_1\, C => 
        \Communications_0/UART_0/tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75499);
    
    HIEFFPLA_INST_0_66101 : AO1A
      port map(A => HIEFFPLA_NET_0_73221, B => 
        HIEFFPLA_NET_0_73231, C => HIEFFPLA_NET_0_73207, Y => 
        HIEFFPLA_NET_0_73209);
    
    \Science_0/ADC_READ_0/cnt[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73290, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73242, Q => 
        \Science_0/ADC_READ_0/cnt[2]_net_1\);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/temp[5]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[5]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72907, Q => 
        \Sensors_0_acc_temp[5]\);
    
    HIEFFPLA_INST_0_59818 : MX2
      port map(A => \Science_0_chan1_data[8]\, B => 
        \Science_0_chan0_data[0]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74503);
    
    HIEFFPLA_INST_0_68485 : NOR3B
      port map(A => HIEFFPLA_NET_0_72639, B => 
        HIEFFPLA_NET_0_72689, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_72640);
    
    HIEFFPLA_INST_0_65522 : NOR3B
      port map(A => HIEFFPLA_NET_0_73352, B => 
        \Science_0/ADC_READ_0/cnt3dn[3]_net_1\, C => 
        \Science_0/ADC_READ_0/cnt3dn[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73353);
    
    \General_Controller_0/status_bits_1[63]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74183, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[63]\);
    
    HIEFFPLA_INST_0_58080 : AND2
      port map(A => \Sensors_0_gyro_y[6]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_74860);
    
    \General_Controller_0/sweep_table_nof_steps[3]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73980, Q => 
        \General_Controller_0/sweep_table_nof_steps[3]_net_1\);
    
    HIEFFPLA_INST_0_60612 : NOR3B
      port map(A => HIEFFPLA_NET_0_74443, B => 
        HIEFFPLA_NET_0_74450, C => HIEFFPLA_NET_0_74725, Y => 
        HIEFFPLA_NET_0_74386);
    
    \Timing_0/s_time[7]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72042, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/s_time[7]_net_1\);
    
    \Science_0/ADC_READ_0/exp_packet_1[42]\ : DFN1E0
      port map(D => \Science_0/ADC_READ_0/data_a[8]_net_1\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[42]\);
    
    HIEFFPLA_INST_0_65698 : NOR2A
      port map(A => HIEFFPLA_NET_0_73309, B => 
        \Science_0/ADC_READ_0/cnt4up[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73306);
    
    HIEFFPLA_INST_0_55183 : AND2
      port map(A => HIEFFPLA_NET_0_75598, B => 
        \Communications_0/UART_0/rx_clk_count[24]_net_1\, Y => 
        HIEFFPLA_NET_0_75566);
    
    HIEFFPLA_INST_0_63144 : NOR3A
      port map(A => HIEFFPLA_NET_0_73937, B => 
        \General_Controller_0/uc_rx_state[2]_net_1\, C => 
        \General_Controller_0/uc_rx_state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73820);
    
    HIEFFPLA_INST_0_70611 : XOR2
      port map(A => \s_clks_net_0[9]\, B => HIEFFPLA_NET_0_72069, 
        Y => HIEFFPLA_NET_0_72065);
    
    HIEFFPLA_INST_0_69901 : NAND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[3]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        Y => HIEFFPLA_NET_0_72272);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[1]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[1]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72808, Q => 
        \Sensors_0_mag_z[1]\);
    
    HIEFFPLA_INST_0_70156 : NAND3A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[5]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[7]_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_write_done\, Y
         => HIEFFPLA_NET_0_72206);
    
    HIEFFPLA_INST_0_57172 : AO1
      port map(A => \Sensors_0_pressure_time[19]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[10]_net_1\, 
        C => HIEFFPLA_NET_0_75010, Y => HIEFFPLA_NET_0_75140);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[0]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72919, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/prev_state[0]_net_1\);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/scl\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_73096, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        ACCE_SCL_c);
    
    HIEFFPLA_INST_0_66973 : AO1C
      port map(A => HIEFFPLA_NET_0_72985, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[1]\, 
        C => HIEFFPLA_NET_0_72993, Y => HIEFFPLA_NET_0_72994);
    
    \General_Controller_0/sweep_table_sample_skip[1]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[1]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[1]_net_1\);
    
    HIEFFPLA_INST_0_61587 : AND3
      port map(A => HIEFFPLA_NET_0_73777, B => 
        HIEFFPLA_NET_0_74173, C => HIEFFPLA_NET_0_73918, Y => 
        HIEFFPLA_NET_0_74178);
    
    \General_Controller_0/sweep_table_write_value[3]\ : DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[3]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[3]_net_1\);
    
    HIEFFPLA_INST_0_61764 : AX1C
      port map(A => 
        \General_Controller_0/sweep_table_sweep_cnt[9]_net_1\, B
         => HIEFFPLA_NET_0_74146, C => 
        \General_Controller_0/sweep_table_sweep_cnt[10]_net_1\, Y
         => HIEFFPLA_NET_0_74143);
    
    \Science_0/DAC_SET_0/cnt[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73217, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Science_0/DAC_SET_0/cnt[2]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/packet_select[8]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_74766, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74760, Q => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\);
    
    HIEFFPLA_INST_0_68531 : AO1
      port map(A => HIEFFPLA_NET_0_72704, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[1]_net_1\, C => 
        HIEFFPLA_NET_0_72632, Y => HIEFFPLA_NET_0_72625);
    
    HIEFFPLA_INST_0_70881 : XA1
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[2]_net_1\, 
        B => HIEFFPLA_NET_0_72762, C => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        Y => HIEFFPLA_NET_0_72006);
    
    HIEFFPLA_INST_0_62198 : AO1
      port map(A => HIEFFPLA_NET_0_73816, B => 
        \General_Controller_0/uc_rx_state_0[4]_net_1\, C => 
        HIEFFPLA_NET_0_74102, Y => HIEFFPLA_NET_0_74032);
    
    HIEFFPLA_INST_0_58654 : AOI1C
      port map(A => HIEFFPLA_NET_0_74650, B => 
        HIEFFPLA_NET_0_74655, C => HIEFFPLA_NET_0_74711, Y => 
        HIEFFPLA_NET_0_74712);
    
    HIEFFPLA_INST_0_66633 : AND3A
      port map(A => HIEFFPLA_NET_0_73077, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        C => HIEFFPLA_NET_0_73038, Y => HIEFFPLA_NET_0_73078);
    
    HIEFFPLA_INST_0_67023 : AO1A
      port map(A => HIEFFPLA_NET_0_72735, B => 
        HIEFFPLA_NET_0_72973, C => HIEFFPLA_NET_0_72982, Y => 
        HIEFFPLA_NET_0_72983);
    
    HIEFFPLA_INST_0_64871 : OR2A
      port map(A => HIEFFPLA_NET_0_73520, B => 
        HIEFFPLA_NET_0_73622, Y => HIEFFPLA_NET_0_73521);
    
    HIEFFPLA_INST_0_64719 : NOR3A
      port map(A => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, B => 
        HIEFFPLA_NET_0_73605, C => HIEFFPLA_NET_0_73563, Y => 
        HIEFFPLA_NET_0_73553);
    
    HIEFFPLA_INST_0_69378 : XOR2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/byte_cnt[0]_net_1\, 
        B => HIEFFPLA_NET_0_72352, Y => HIEFFPLA_NET_0_72404);
    
    HIEFFPLA_INST_0_58523 : NOR3B
      port map(A => HIEFFPLA_NET_0_74738, B => 
        HIEFFPLA_NET_0_74730, C => HIEFFPLA_NET_0_74740, Y => 
        HIEFFPLA_NET_0_74743);
    
    HIEFFPLA_INST_0_62407 : OR3A
      port map(A => HIEFFPLA_NET_0_73905, B => 
        HIEFFPLA_NET_0_73776, C => 
        \General_Controller_0/uc_rx_state_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73989);
    
    HIEFFPLA_INST_0_68418 : NOR2A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_data_out[0]\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72655);
    
    HIEFFPLA_INST_0_67973 : AND3C
      port map(A => HIEFFPLA_NET_0_72739, B => 
        \Sensors_0/Accelerometer_0/state_0[8]\, C => 
        HIEFFPLA_NET_0_72912, Y => HIEFFPLA_NET_0_72764);
    
    HIEFFPLA_INST_0_64584 : AND3C
      port map(A => \General_Controller_0/uc_tx_state[6]_net_1\, 
        B => \General_Controller_0/uc_tx_state[7]_net_1\, C => 
        \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73596);
    
    \Science_0/DAC_SET_0/vector[8]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73188, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[8]_net_1\);
    
    HIEFFPLA_INST_0_60233 : MX2
      port map(A => HIEFFPLA_NET_0_74565, B => 
        HIEFFPLA_NET_0_74416, S => HIEFFPLA_NET_0_74340, Y => 
        HIEFFPLA_NET_0_74443);
    
    HIEFFPLA_INST_0_68594 : AO1
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/GYRO_SCL_c_0\, C => 
        HIEFFPLA_NET_0_72699, Y => HIEFFPLA_NET_0_72610);
    
    HIEFFPLA_INST_0_55150 : XA1B
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[25]_net_1\, B => 
        HIEFFPLA_NET_0_75577, C => HIEFFPLA_NET_0_75567, Y => 
        HIEFFPLA_NET_0_75574);
    
    \Timekeeper_0/microseconds[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72132, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[5]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72218, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[1]_net_1\);
    
    HIEFFPLA_INST_0_70337 : AOI1D
      port map(A => General_Controller_0_st_ren1, B => 
        \SweepTable_0/WEBP\, C => 
        \General_Controller_0_st_raddr_1[1]\, Y => 
        \TableSelect_0_RADDR[1]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[12]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72553, Q => 
        \Sensors_0_gyro_x[12]\);
    
    HIEFFPLA_INST_0_58186 : AO1
      port map(A => \Science_0_exp_packet_0[58]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_75126, Y => HIEFFPLA_NET_0_74834);
    
    HIEFFPLA_INST_0_59979 : MX2
      port map(A => \Science_0_chan0_data[4]\, B => 
        \Science_0_chan0_data[8]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74479);
    
    HIEFFPLA_INST_0_55386 : NAND2B
      port map(A => HIEFFPLA_NET_0_75515, B => 
        HIEFFPLA_NET_0_75527, Y => HIEFFPLA_NET_0_75524);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[1]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75266, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[1]\\\\\);
    
    HIEFFPLA_INST_0_69967 : AOI1D
      port map(A => HIEFFPLA_NET_0_72228, B => 
        HIEFFPLA_NET_0_72231, C => HIEFFPLA_NET_0_72253, Y => 
        HIEFFPLA_NET_0_72258);
    
    HIEFFPLA_INST_0_66281 : NAND2
      port map(A => HIEFFPLA_NET_0_73175, B => 
        \Science_0/SET_LP_GAIN_0/state[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73157);
    
    \Communications_0/UART_0/rx_byte[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75380, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75610, Q => 
        \Communications_0/UART_0/rx_byte[2]_net_1\);
    
    \Science_0/ADC_READ_0/cnt2dn[1]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73375, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73424, Q => 
        \Science_0/ADC_READ_0/cnt2dn[1]_net_1\);
    
    HIEFFPLA_INST_0_64377 : MX2
      port map(A => HIEFFPLA_NET_0_73712, B => 
        HIEFFPLA_NET_0_73704, S => HIEFFPLA_NET_0_73593, Y => 
        HIEFFPLA_NET_0_73632);
    
    HIEFFPLA_INST_0_58281 : AO1
      port map(A => \Sensors_0_acc_x[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74812, Y => HIEFFPLA_NET_0_74813);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRY[4]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75300, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[4]\\\\\);
    
    HIEFFPLA_INST_0_62764 : OA1A
      port map(A => HIEFFPLA_NET_0_73784, B => 
        HIEFFPLA_NET_0_74125, C => HIEFFPLA_NET_0_73918, Y => 
        HIEFFPLA_NET_0_73911);
    
    HIEFFPLA_INST_0_64110 : OR2A
      port map(A => HIEFFPLA_NET_0_73579, B => 
        \General_Controller_0/constant_bias_voltage_0[10]_net_1\, 
        Y => HIEFFPLA_NET_0_73669);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[11]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[3]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72281, Q => \Sensors_0_pressure_raw[11]\);
    
    HIEFFPLA_INST_0_65410 : AND2B
      port map(A => \Science_0/ADC_READ_0/cnt2dn[0]_net_1\, B => 
        \Science_0/ADC_READ_0/cnt2dn[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73384);
    
    HIEFFPLA_INST_0_59144 : AO1
      port map(A => HIEFFPLA_NET_0_74596, B => 
        \GS_Readout_0/state[5]_net_1\, C => HIEFFPLA_NET_0_74600, 
        Y => HIEFFPLA_NET_0_74601);
    
    HIEFFPLA_INST_0_61874 : NOR3A
      port map(A => HIEFFPLA_NET_0_74115, B => 
        HIEFFPLA_NET_0_73889, C => 
        \General_Controller_0/uc_rx_byte[2]_net_1\, Y => 
        HIEFFPLA_NET_0_74111);
    
    HIEFFPLA_INST_0_60480 : MX2
      port map(A => \Science_0_chan7_data[2]\, B => 
        \Science_0_chan7_data[6]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74409);
    
    HIEFFPLA_INST_0_56395 : AX1C
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, B
         => HIEFFPLA_NET_0_75371, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\, Y
         => HIEFFPLA_NET_0_75291);
    
    HIEFFPLA_INST_0_70878 : MX2A
      port map(A => HIEFFPLA_NET_0_72007, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0_num_bytes[2]\, S
         => \Sensors_0/Gyro_0/I2C_Master_0/state[7]_net_1\, Y => 
        HIEFFPLA_NET_0_72686);
    
    \General_Controller_0/uc_tx_substate[0]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_73551, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_tx_substate[0]_net_1\);
    
    \Timing_0/m_time[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72067, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \Timing_0/m_time[0]_net_1\);
    
    \Timekeeper_0/microseconds[12]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72148, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[12]\);
    
    HIEFFPLA_INST_0_57651 : AO1B
      port map(A => \Sensors_0_gyro_y[10]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74980, Y => HIEFFPLA_NET_0_74981);
    
    \GYRO_SCL_pad/U0/U0\ : IOPAD_TRI
      port map(D => \GYRO_SCL_pad/U0/NET1\, E => 
        \GYRO_SCL_pad/U0/NET2\, PAD => GYRO_SCL);
    
    HIEFFPLA_INST_0_62060 : NAND2A
      port map(A => HIEFFPLA_NET_0_74062, B => 
        HIEFFPLA_NET_0_73943, Y => HIEFFPLA_NET_0_74060);
    
    HIEFFPLA_INST_0_57860 : AOI1
      port map(A => \Sensors_0_acc_time[21]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74922, Y => HIEFFPLA_NET_0_74923);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/acc_time[17]\ : 
        DFN1E1
      port map(D => \Timekeeper_0_microseconds[17]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72920, Q => 
        \Sensors_0_acc_time[17]\);
    
    HIEFFPLA_INST_0_58888 : AND3
      port map(A => HIEFFPLA_NET_0_74694, B => 
        HIEFFPLA_NET_0_74510, C => HIEFFPLA_NET_0_74386, Y => 
        HIEFFPLA_NET_0_74665);
    
    HIEFFPLA_INST_0_69744 : AO1A
      port map(A => PRESSURE_SCL_c, B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[4]_net_1\, 
        C => HIEFFPLA_NET_0_72422, Y => HIEFFPLA_NET_0_72318);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[20]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72282, Q => 
        \Sensors_0_pressure_temp_raw[20]\);
    
    HIEFFPLA_INST_0_68629 : NAND3C
      port map(A => HIEFFPLA_NET_0_72664, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[0]_net_1\, C
         => \Sensors_0/Gyro_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_72602);
    
    HIEFFPLA_INST_0_63025 : AO1
      port map(A => HIEFFPLA_NET_0_73896, B => 
        HIEFFPLA_NET_0_73796, C => HIEFFPLA_NET_0_73838, Y => 
        HIEFFPLA_NET_0_73845);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/data_out[4]\ : 
        DFN0E1C1
      port map(D => ACCE_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73120, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[4]\);
    
    HIEFFPLA_INST_0_70547 : AND2
      port map(A => \Timing_0/m_count[5]_net_1\, B => 
        \Timing_0/m_count[2]_net_1\, Y => HIEFFPLA_NET_0_72084);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_z[2]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72808, Q => 
        \Sensors_0_mag_z[2]\);
    
    HIEFFPLA_INST_0_67442 : NOR3B
      port map(A => HIEFFPLA_NET_0_72904, B => 
        HIEFFPLA_NET_0_72905, C => HIEFFPLA_NET_0_72876, Y => 
        HIEFFPLA_NET_0_72878);
    
    HIEFFPLA_INST_0_56412 : MX2
      port map(A => \FMC_DA_c[1]\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[1]\\\\\, S => 
        \Data_Saving_0/FPGA_Buffer_0/DVLDI\, Y => 
        HIEFFPLA_NET_0_75286);
    
    HIEFFPLA_INST_0_55042 : NOR3B
      port map(A => HIEFFPLA_NET_0_75563, B => 
        HIEFFPLA_NET_0_75604, C => 
        \Communications_0/UART_0/rx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75606);
    
    \General_Controller_0/sweep_table_probe_id[4]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[4]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73924, Q => 
        \General_Controller_0/sweep_table_probe_id[4]_net_1\);
    
    HIEFFPLA_INST_0_57664 : AOI1
      port map(A => \Science_0_exp_packet_0[35]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_74976, Y => HIEFFPLA_NET_0_74977);
    
    \General_Controller_0/uc_tx_state[0]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_73575, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73595, Q => 
        \General_Controller_0/uc_tx_state[0]_net_1\);
    
    HIEFFPLA_INST_0_67809 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        B => HIEFFPLA_NET_0_72737, C => HIEFFPLA_NET_0_72799, Y
         => HIEFFPLA_NET_0_72796);
    
    HIEFFPLA_INST_0_66622 : AOI1A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        C => HIEFFPLA_NET_0_73145, Y => HIEFFPLA_NET_0_73080);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/isSetup\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72969, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/isSetup_net_1\);
    
    \Science_0/ADC_READ_0/cnt4dn[0]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73318, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73422, Q => 
        \Science_0/ADC_READ_0/cnt4dn[0]_net_1\);
    
    HIEFFPLA_INST_0_65779 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt[5]_net_1\, B => 
        HIEFFPLA_NET_0_73293, C => 
        \Science_0/ADC_READ_0/cnt[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73281);
    
    HIEFFPLA_INST_0_55453 : AND2B
      port map(A => HIEFFPLA_NET_0_75502, B => 
        \Communications_0/UART_0/tx_count[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75508);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/temp[5]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[5]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72555, Q => 
        \Sensors_0_gyro_temp[5]\);
    
    HIEFFPLA_INST_0_58195 : AO1
      port map(A => \Science_0_exp_packet_0[61]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_75124, Y => HIEFFPLA_NET_0_74832);
    
    HIEFFPLA_INST_0_54946 : AND3
      port map(A => \ClockDivs_0/cnt_800kHz[0]_net_1\, B => 
        \ClockDivs_0/cnt_800kHz[1]_net_1\, C => 
        \ClockDivs_0/cnt_800kHz[2]_net_1\, Y => 
        HIEFFPLA_NET_0_75632);
    
    \General_Controller_0/st_wdata[10]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[10]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[10]\);
    
    \General_Controller_0/status_bits_1[40]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74206, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[40]\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRY[0]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75307, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[0]\\\\\);
    
    \Communications_0/UART_1/rx_byte[5]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75378, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75491, Q => 
        \Communications_0/UART_1/rx_byte[5]_net_1\);
    
    \Science_0/ADC_READ_0/chan3_data[0]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_a[6]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan3_data[0]\);
    
    HIEFFPLA_INST_0_60444 : MX2
      port map(A => HIEFFPLA_NET_0_74511, B => 
        HIEFFPLA_NET_0_74438, S => HIEFFPLA_NET_0_74342, Y => 
        HIEFFPLA_NET_0_74413);
    
    HIEFFPLA_INST_0_57491 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[11]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_75030, Y => HIEFFPLA_NET_0_75031);
    
    HIEFFPLA_INST_0_69067 : NAND2
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        B => \Sensors_0/Gyro_0/I2C_Master_0_data_out_rdy\, Y => 
        HIEFFPLA_NET_0_72479);
    
    HIEFFPLA_INST_0_62487 : NOR3B
      port map(A => HIEFFPLA_NET_0_73900, B => 
        HIEFFPLA_NET_0_73906, C => 
        \General_Controller_0/uc_rx_state_0[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73972);
    
    HIEFFPLA_INST_0_68898 : NOR3A
      port map(A => HIEFFPLA_NET_0_72525, B => 
        HIEFFPLA_NET_0_72487, C => HIEFFPLA_NET_0_72526, Y => 
        HIEFFPLA_NET_0_72527);
    
    HIEFFPLA_INST_0_68598 : AO1A
      port map(A => HIEFFPLA_NET_0_72705, B => 
        HIEFFPLA_NET_0_72620, C => HIEFFPLA_NET_0_72600, Y => 
        HIEFFPLA_NET_0_72609);
    
    HIEFFPLA_INST_0_56297 : AX1
      port map(A => HIEFFPLA_NET_0_75370, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, C
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, 
        Y => HIEFFPLA_NET_0_75315);
    
    HIEFFPLA_INST_0_61802 : OR3A
      port map(A => HIEFFPLA_NET_0_73780, B => 
        HIEFFPLA_NET_0_74124, C => HIEFFPLA_NET_0_73786, Y => 
        HIEFFPLA_NET_0_74126);
    
    \Communications_0/UART_1/rx_clk_count[28]\ : DFN1E0C1
      port map(D => HIEFFPLA_NET_0_75459, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75443, Q => 
        \Communications_0/UART_1/rx_clk_count[28]_net_1\);
    
    HIEFFPLA_INST_0_65072 : AO1D
      port map(A => HIEFFPLA_NET_0_73479, B => 
        \Pressure_Signal_Debounce_0/state[0]_net_1\, C => 
        HIEFFPLA_NET_0_73475, Y => HIEFFPLA_NET_0_73476);
    
    HIEFFPLA_INST_0_64575 : NAND2B
      port map(A => \General_Controller_0/uc_tx_state[0]_net_1\, 
        B => \General_Controller_0/uc_tx_state[6]_net_1\, Y => 
        HIEFFPLA_NET_0_73598);
    
    HIEFFPLA_INST_0_55678 : OA1A
      port map(A => HIEFFPLA_NET_0_75451, B => 
        \Communications_0/UART_1/rx_count[2]_net_1\, C => 
        \Communications_0/UART_1/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75448);
    
    HIEFFPLA_INST_0_69060 : NOR3A
      port map(A => HIEFFPLA_NET_0_72483, B => 
        HIEFFPLA_NET_0_72548, C => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[6]_net_1\, 
        Y => HIEFFPLA_NET_0_72482);
    
    HIEFFPLA_INST_0_63620 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[14]_net_1\, 
        B => 
        \General_Controller_0/sweep_table_sample_skip[14]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73739);
    
    \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[3]\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_72685, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72618, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/byte_cnt[3]_net_1\);
    
    HIEFFPLA_INST_0_56335 : XOR2
      port map(A => HIEFFPLA_NET_0_75331, B => 
        HIEFFPLA_NET_0_75294, Y => HIEFFPLA_NET_0_75307);
    
    \Timing_0/m_time[7]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_72071, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => \m_time[7]\);
    
    HIEFFPLA_INST_0_59973 : MX2
      port map(A => \Sensors_0_pressure_temp_raw[15]\, B => 
        \Sensors_0_pressure_temp_raw[19]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74480);
    
    HIEFFPLA_INST_0_66797 : AO1
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        B => ACCE_SCL_c, C => HIEFFPLA_NET_0_73051, Y => 
        HIEFFPLA_NET_0_73033);
    
    \General_Controller_0/st_wdata[0]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/sweep_table_write_value[0]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73802, Q => 
        \General_Controller_0_st_wdata[0]\);
    
    HIEFFPLA_INST_0_58616 : AND3
      port map(A => HIEFFPLA_NET_0_74724, B => 
        HIEFFPLA_NET_0_74723, C => HIEFFPLA_NET_0_74722, Y => 
        HIEFFPLA_NET_0_74719);
    
    HIEFFPLA_INST_0_58078 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[22]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[10]_net_1\, 
        C => HIEFFPLA_NET_0_74860, Y => HIEFFPLA_NET_0_74861);
    
    AFLSDF_INV_7 : INV
      port map(A => CLKINT_1_Y, Y => \AFLSDF_INV_7\);
    
    HIEFFPLA_INST_0_63638 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[9]_net_1\, B
         => 
        \General_Controller_0/sweep_table_samples_per_point[9]_net_1\, 
        S => \General_Controller_0/uc_tx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73736);
    
    HIEFFPLA_INST_0_71209 : AXOI1
      port map(A => HIEFFPLA_NET_0_75453, B => 
        \Communications_0/UART_1/rx_count[0]_net_1\, C => 
        HIEFFPLA_NET_0_75442, Y => HIEFFPLA_NET_0_71973);
    
    \Science_0/ADC_READ_0/chan5_data[5]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[5]\);
    
    HIEFFPLA_INST_0_68331 : NOR3A
      port map(A => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, B => 
        HIEFFPLA_NET_0_72676, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[2]_net_1\, Y => 
        HIEFFPLA_NET_0_72680);
    
    HIEFFPLA_INST_0_58102 : AND2
      port map(A => \ch3_data_net_0[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_74855);
    
    HIEFFPLA_INST_0_56549 : NAND2
      port map(A => HIEFFPLA_NET_0_75255, B => 
        \Data_Saving_0/Interrupt_Generator_0/counter[8]_net_1\, Y
         => HIEFFPLA_NET_0_75243);
    
    \Communications_0/UART_1/rx_state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75435, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/rx_state[1]_net_1\);
    
    HIEFFPLA_INST_0_65655 : XA1
      port map(A => HIEFFPLA_NET_0_73324, B => 
        \Science_0/ADC_READ_0/cnt4dn[2]_net_1\, C => 
        HIEFFPLA_NET_0_73274, Y => HIEFFPLA_NET_0_73316);
    
    HIEFFPLA_INST_0_66196 : AOI1
      port map(A => \Science_0/SET_LP_GAIN_0/state[7]_net_1\, B
         => \Science_0/ADC_READ_0_G1[1]\, C => 
        HIEFFPLA_NET_0_73180, Y => HIEFFPLA_NET_0_73181);
    
    HIEFFPLA_INST_0_63854 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_read_value[5]_net_1\, B
         => 
        \General_Controller_0/sweep_table_sample_skip[5]_net_1\, 
        S => \General_Controller_0/uc_tx_state[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73700);
    
    HIEFFPLA_INST_0_64624 : NOR3B
      port map(A => HIEFFPLA_NET_0_73609, B => 
        HIEFFPLA_NET_0_73920, C => HIEFFPLA_NET_0_73978, Y => 
        HIEFFPLA_NET_0_73583);
    
    \General_Controller_0/sweep_table_samples_per_point[13]\ : 
        DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[5]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[13]_net_1\);
    
    \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_74762, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1E1C0_data_out[0]\\\\/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75287, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \FMC_DA_c[0]\);
    
    HIEFFPLA_INST_0_69565 : AND3
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_1_net_1\, 
        C => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/sda_cl_2_net_1\, 
        Y => sda_cl_1_RNIGPAD);
    
    HIEFFPLA_INST_0_61556 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[62]\, B => 
        \Timekeeper_0_milliseconds[22]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74184);
    
    \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_73030, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[5]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRY[6]\\\\\ : DFN1C0
      port map(D => HIEFFPLA_NET_0_75305, CLK => CLKINT_0_Y_0, 
        CLR => \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRY[6]\\\\\);
    
    HIEFFPLA_INST_0_69597 : AO1A
      port map(A => CLKINT_1_Y, B => HIEFFPLA_NET_0_72347, C => 
        HIEFFPLA_NET_0_72353, Y => HIEFFPLA_NET_0_72354);
    
    HIEFFPLA_INST_0_67713 : NOR3B
      port map(A => HIEFFPLA_NET_0_72846, B => 
        HIEFFPLA_NET_0_72845, C => HIEFFPLA_NET_0_72937, Y => 
        HIEFFPLA_NET_0_72817);
    
    HIEFFPLA_INST_0_65832 : NOR2A
      port map(A => \Science_0/ADC_READ_0/newflag_net_1\, B => 
        General_Controller_0_en_science_packets, Y => 
        HIEFFPLA_NET_0_73273);
    
    \General_Controller_0/uc_tx_substate[2]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73549, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/uc_tx_substate[2]_net_1\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1E1C0_data_out[7]\\\\/U1\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75280, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \FMC_DA_c[7]\);
    
    \Data_Saving_0/Packet_Saver_0/data_out[27]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75216, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[27]\);
    
    \Science_0/ADC_READ_0/chan6_data[4]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan6_data[4]\);
    
    \Science_0/ADC_READ_0/chan0_data[4]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73418, Q => \Science_0_chan0_data[4]\);
    
    HIEFFPLA_INST_0_60869 : NAND3C
      port map(A => \General_Controller_0/command[3]_net_1\, B
         => \General_Controller_0/command[7]_net_1\, C => 
        \General_Controller_0/ext_rx_state_i_0[1]\, Y => 
        HIEFFPLA_NET_0_74335);
    
    HIEFFPLA_INST_0_54952 : XOR2
      port map(A => \ClockDivs_0/cnt_800kHz[0]_net_1\, B => 
        \ClockDivs_0/cnt_800kHz[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75630);
    
    HIEFFPLA_INST_0_62506 : AND3
      port map(A => HIEFFPLA_NET_0_74026, B => 
        HIEFFPLA_NET_0_74110, C => HIEFFPLA_NET_0_73805, Y => 
        HIEFFPLA_NET_0_73968);
    
    HIEFFPLA_INST_0_55524 : AND3A
      port map(A => HIEFFPLA_NET_0_75473, B => 
        \Communications_0/UART_1/rx_clk_count[24]_net_1\, C => 
        HIEFFPLA_NET_0_75474, Y => HIEFFPLA_NET_0_75488);
    
    \Data_Saving_0/FPGA_Buffer_0/_RAM4K9_QXI[7]_\ : RAM4K9
      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[7]\\\\\, 
        ADDRA6 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[6]\\\\\, 
        ADDRA5 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\, 
        ADDRA4 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, 
        ADDRA3 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, 
        ADDRA2 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[2]\\\\\, 
        ADDRA1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[1]\\\\\, 
        ADDRA0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[0]\\\\\, 
        ADDRB11 => AFLSDF_GND, ADDRB10 => \GND\, ADDRB9 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\, 
        ADDRB8 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, 
        ADDRB7 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[7]\\\\\, 
        ADDRB6 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, 
        ADDRB5 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\, 
        ADDRB4 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, 
        ADDRB3 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, 
        ADDRB2 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[2]\\\\\, 
        ADDRB1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[1]\\\\\, 
        ADDRB0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[0]\\\\\, 
        DINA8 => \GND\, DINA7 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[31]\, DINA6 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[30]\, DINA5 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[23]\, DINA4 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[22]\, DINA3 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[15]\, DINA2 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[14]\, DINA1 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[7]\, DINA0 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[6]\, DINB8 => 
        \GND\, DINB7 => \GND\, DINB6 => \GND\, DINB5 => \GND\, 
        DINB4 => \GND\, DINB3 => \GND\, DINB2 => \GND\, DINB1 => 
        \GND\, DINB0 => \GND\, WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, 
        WIDTHB0 => \VCC\, WIDTHB1 => \GND\, PIPEA => \GND\, PIPEB
         => \GND\, WMODEA => \GND\, WMODEB => \GND\, BLKA => 
        \Data_Saving_0/FPGA_Buffer_0/MEMWENEG\, BLKB => 
        \AFLSDF_INV_3\, WENA => \GND\, WENB => \VCC\, CLKA => 
        CLKINT_0_Y_0, CLKB => CLKINT_2_Y, RESET => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, DOUTA8 => 
        OPEN, DOUTA7 => OPEN, DOUTA6 => OPEN, DOUTA5 => OPEN, 
        DOUTA4 => OPEN, DOUTA3 => OPEN, DOUTA2 => OPEN, DOUTA1
         => OPEN, DOUTA0 => OPEN, DOUTB8 => OPEN, DOUTB7 => OPEN, 
        DOUTB6 => OPEN, DOUTB5 => OPEN, DOUTB4 => OPEN, DOUTB3
         => OPEN, DOUTB2 => OPEN, DOUTB1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[7]\\\\\, DOUTB0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[6]\\\\\);
    
    \Science_0/ADC_READ_0/chan5_data[10]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[16]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan5_data[10]\);
    
    HIEFFPLA_INST_0_57152 : AND2
      port map(A => \Sensors_0_gyro_y[15]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, Y
         => HIEFFPLA_NET_0_75153);
    
    \Science_0/ADC_READ_0/data_b[12]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_b[11]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        \Science_0/ADC_READ_0/state_0[1]_net_1\, Q => 
        \Science_0/ADC_READ_0/data_b[12]_net_1\);
    
    HIEFFPLA_INST_0_66045 : NAND2B
      port map(A => \Science_0/DAC_SET_0/state[4]_net_1\, B => 
        \Science_0/DAC_SET_0/state[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73227);
    
    HIEFFPLA_INST_0_56476 : XOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[2]\\\\\, B => 
        HIEFFPLA_NET_0_75323, C => HIEFFPLA_NET_0_75322, Y => 
        HIEFFPLA_NET_0_75270);
    
    HIEFFPLA_INST_0_65270 : NOR3A
      port map(A => HIEFFPLA_NET_0_73431, B => 
        \Sensors_0_pressure_raw[7]\, C => 
        \Sensors_0_pressure_raw[4]\, Y => HIEFFPLA_NET_0_73429);
    
    HIEFFPLA_INST_0_65225 : AND2
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[6]_net_1\, 
        B => \Pressure_Signal_Debounce_0/ms_cnt[7]_net_1\, Y => 
        HIEFFPLA_NET_0_73441);
    
    HIEFFPLA_INST_0_55582 : NOR3A
      port map(A => HIEFFPLA_NET_0_75471, B => 
        \Communications_0/UART_1/rx_state[0]_net_1\, C => 
        \Communications_0/UART_1/rx_clk_count[23]_net_1\, Y => 
        HIEFFPLA_NET_0_75474);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72336, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[3]_net_1\);
    
    HIEFFPLA_INST_0_66874 : OA1C
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_we\, 
        C => HIEFFPLA_NET_0_73046, Y => HIEFFPLA_NET_0_73015);
    
    \Sensors_0/Gyro_0/I2C_Master_0/sda_cl\ : DFN0C1
      port map(D => HIEFFPLA_NET_0_72635, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/sda_cl_net_1\);
    
    HIEFFPLA_INST_0_68093 : AOI1A
      port map(A => HIEFFPLA_NET_0_72911, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[3]_net_1\, 
        C => HIEFFPLA_NET_0_72926, Y => HIEFFPLA_NET_0_72731);
    
    HIEFFPLA_INST_0_63436 : MX2
      port map(A => HIEFFPLA_NET_0_73755, B => 
        HIEFFPLA_NET_0_73689, S => HIEFFPLA_NET_0_73608, Y => 
        HIEFFPLA_NET_0_73763);
    
    \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/temp[3]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72907, Q => 
        \Sensors_0_acc_temp[3]\);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[8]\ : DFN0P1
      port map(D => HIEFFPLA_NET_0_72332, CLK => 
        ClockDivs_0_clk_800kHz, PRE => CLKINT_1_Y, Q => 
        \Sensors_0/Pressure_Sensor_0/state[8]\);
    
    HIEFFPLA_INST_0_68901 : NOR3A
      port map(A => General_Controller_0_en_sensors, B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/state_i_0[4]\, C
         => \Sensors_0/Gyro_0/L3GD20H_Interface_0/isSetup_net_1\, 
        Y => HIEFFPLA_NET_0_72526);
    
    HIEFFPLA_INST_0_64799 : AO1
      port map(A => 
        \General_Controller_0/uc_tx_substate[2]_net_1\, B => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, C => 
        HIEFFPLA_NET_0_73557, Y => HIEFFPLA_NET_0_73540);
    
    \Communications_0/UART_1/recv[7]\ : DFN1E1C1
      port map(D => \Communications_0/UART_1/rx_byte[7]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_75441, Q => \Communications_0_uc_recv[7]\);
    
    HIEFFPLA_INST_0_58217 : AO1
      port map(A => \Sensors_0_mag_y[9]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[11]_net_1\, 
        C => HIEFFPLA_NET_0_75097, Y => HIEFFPLA_NET_0_74825);
    
    HIEFFPLA_INST_0_58290 : AO1
      port map(A => \Science_0_exp_packet_0[40]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_75088, Y => HIEFFPLA_NET_0_74810);
    
    HIEFFPLA_INST_0_61317 : XA1C
      port map(A => HIEFFPLA_NET_0_74261, B => 
        \General_Controller_0/state_seconds[8]_net_1\, C => 
        HIEFFPLA_NET_0_74217, Y => HIEFFPLA_NET_0_74219);
    
    \Timekeeper_0/microseconds[16]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72144, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72092, Q => 
        \Timekeeper_0_microseconds[16]\);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[4]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[4]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72503, Q => 
        \Sensors_0_gyro_x[4]\);
    
    HIEFFPLA_INST_0_60645 : MX2
      port map(A => \Science_0_chan6_data[5]\, B => 
        \Science_0_chan6_data[9]\, S => 
        \GS_Readout_0/subState[0]_net_1\, Y => 
        HIEFFPLA_NET_0_74381);
    
    HIEFFPLA_INST_0_68139 : NAND3C
      port map(A => HIEFFPLA_NET_0_72730, B => 
        HIEFFPLA_NET_0_72733, C => HIEFFPLA_NET_0_72721, Y => 
        HIEFFPLA_NET_0_72725);
    
    HIEFFPLA_INST_0_61735 : XA1B
      port map(A => 
        \General_Controller_0/sweep_table_read_wait[31]_net_1\, B
         => HIEFFPLA_NET_0_73815, C => HIEFFPLA_NET_0_73977, Y
         => HIEFFPLA_NET_0_74151);
    
    HIEFFPLA_INST_0_70729 : AND2
      port map(A => HIEFFPLA_NET_0_72030, B => 
        \Timing_0/m_count[6]_net_1\, Y => HIEFFPLA_NET_0_72029);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/data_out[4]\ : 
        DFN0E1C1
      port map(D => PRESSURE_SDA_in, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72398, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[4]\);
    
    HIEFFPLA_INST_0_64639 : NOR3B
      port map(A => HIEFFPLA_NET_0_73578, B => 
        \General_Controller_0/uc_tx_state[7]_net_1\, C => 
        HIEFFPLA_NET_0_74323, Y => HIEFFPLA_NET_0_73579);
    
    HIEFFPLA_INST_0_66449 : NOR3B
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[0]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[2]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73118);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/data_out_1[3]\ : 
        DFN1E0C1
      port map(D => HIEFFPLA_NET_0_72285, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72270, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0_data_out[3]\);
    
    \Communications_0/UART_1/rx_count[2]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_75448, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_75442, Q => 
        \Communications_0/UART_1/rx_count[2]_net_1\);
    
    HIEFFPLA_INST_0_66640 : AND3C
      port map(A => HIEFFPLA_NET_0_73075, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[2]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/byte_cnt[3]_net_1\, 
        Y => HIEFFPLA_NET_0_73076);
    
    HIEFFPLA_INST_0_60847 : NOR3B
      port map(A => \GS_Readout_0/state[6]_net_1\, B => 
        HIEFFPLA_NET_0_74344, C => Communications_0_ext_tx_rdy, Y
         => HIEFFPLA_NET_0_74345);
    
    HIEFFPLA_INST_0_57404 : AO1
      port map(A => \Science_0_exp_packet_0[3]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_74850, Y => HIEFFPLA_NET_0_75055);
    
    HIEFFPLA_INST_0_56786 : MX2
      port map(A => HIEFFPLA_NET_0_75173, B => 
        HIEFFPLA_NET_0_75031, S => HIEFFPLA_NET_0_74755, Y => 
        HIEFFPLA_NET_0_75210);
    
    HIEFFPLA_INST_0_54955 : XOR2
      port map(A => HIEFFPLA_NET_0_75632, B => 
        \ClockDivs_0/cnt_800kHz[3]_net_1\, Y => 
        HIEFFPLA_NET_0_75628);
    
    HIEFFPLA_INST_0_65362 : AX1C
      port map(A => \Science_0/ADC_READ_0/cnt1dn[3]_net_1\, B => 
        HIEFFPLA_NET_0_73410, C => 
        \Science_0/ADC_READ_0/cnt1dn[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73400);
    
    \UC_UART_RX_pad/U0/U0\ : IOPAD_TRI
      port map(D => \UC_UART_RX_pad/U0/NET1\, E => 
        \UC_UART_RX_pad/U0/NET2\, PAD => UC_UART_RX);
    
    HIEFFPLA_INST_0_67338 : AND3C
      port map(A => HIEFFPLA_NET_0_72898, B => 
        HIEFFPLA_NET_0_72892, C => HIEFFPLA_NET_0_72927, Y => 
        HIEFFPLA_NET_0_72904);
    
    HIEFFPLA_INST_0_66465 : AND2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_repeat_start\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73113);
    
    HIEFFPLA_INST_0_61017 : NOR3B
      port map(A => HIEFFPLA_NET_0_74253, B => 
        HIEFFPLA_NET_0_74296, C => 
        \General_Controller_0/state_seconds[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74294);
    
    HIEFFPLA_INST_0_55098 : NOR3A
      port map(A => 
        \Communications_0/UART_0/rx_clk_count[24]_net_1\, B => 
        HIEFFPLA_NET_0_75590, C => 
        \Communications_0/UART_0/rx_clk_count[27]_net_1\, Y => 
        HIEFFPLA_NET_0_75591);
    
    HIEFFPLA_INST_0_58232 : AO1
      port map(A => \Sensors_0_mag_x[5]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[11]_net_1\, C
         => HIEFFPLA_NET_0_75130, Y => HIEFFPLA_NET_0_74823);
    
    \General_Controller_0/sweep_table_samples_per_point[4]\ : 
        DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[4]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74033, Q => 
        \General_Controller_0/sweep_table_samples_per_point[4]_net_1\);
    
    \General_Controller_0/uc_rx_byte[2]\ : DFN1E1
      port map(D => \Communications_0_uc_recv[2]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74031, Q => 
        \General_Controller_0/uc_rx_byte[2]_net_1\);
    
    HIEFFPLA_INST_0_59288 : NOR2A
      port map(A => HIEFFPLA_NET_0_74493, B => 
        HIEFFPLA_NET_0_74725, Y => HIEFFPLA_NET_0_74574);
    
    HIEFFPLA_INST_0_58836 : AND2
      port map(A => HIEFFPLA_NET_0_74645, B => 
        HIEFFPLA_NET_0_74459, Y => HIEFFPLA_NET_0_74677);
    
    \Sensors_0/Gyro_0/I2C_Master_0/data_out[6]\ : DFN0E1C1
      port map(D => GYRO_SDA_in, CLK => ClockDivs_0_clk_800kHz, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72675, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0_data_out[6]\);
    
    HIEFFPLA_INST_0_61500 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[55]\, B => 
        \Timekeeper_0_milliseconds[15]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74191);
    
    HIEFFPLA_INST_0_62586 : OR3A
      port map(A => \General_Controller_0/uc_rx_state[0]_net_1\, 
        B => HIEFFPLA_NET_0_74072, C => 
        \General_Controller_0/uc_rx_state[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73951);
    
    HIEFFPLA_INST_0_59326 : AND3B
      port map(A => HIEFFPLA_NET_0_74433, B => 
        HIEFFPLA_NET_0_74725, C => HIEFFPLA_NET_0_74564, Y => 
        HIEFFPLA_NET_0_74568);
    
    HIEFFPLA_INST_0_58855 : NOR3B
      port map(A => HIEFFPLA_NET_0_74371, B => 
        \GS_Readout_0/state[3]_net_1\, C => HIEFFPLA_NET_0_74474, 
        Y => HIEFFPLA_NET_0_74673);
    
    HIEFFPLA_INST_0_70088 : AO1E
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[8]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/subState[6]_net_1\, 
        C => HIEFFPLA_NET_0_72275, Y => HIEFFPLA_NET_0_72224);
    
    HIEFFPLA_INST_0_63176 : NOR3A
      port map(A => HIEFFPLA_NET_0_73972, B => 
        HIEFFPLA_NET_0_74154, C => HIEFFPLA_NET_0_73784, Y => 
        HIEFFPLA_NET_0_73815);
    
    HIEFFPLA_INST_0_61195 : NOR3A
      port map(A => HIEFFPLA_NET_0_74252, B => 
        \General_Controller_0/state_seconds[5]_net_1\, C => 
        \General_Controller_0/state_seconds[4]_net_1\, Y => 
        HIEFFPLA_NET_0_74253);
    
    \Sensors_0/Gyro_0/I2C_Master_0/next_state[0]\ : DFN0E0
      port map(D => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[4]_net_1\, CLK => 
        ClockDivs_0_clk_800kHz, E => HIEFFPLA_NET_0_72617, Q => 
        \Sensors_0/Gyro_0/I2C_Master_0/next_state[0]_net_1\);
    
    HIEFFPLA_INST_0_56535 : XOR2
      port map(A => HIEFFPLA_NET_0_75254, B => 
        \Data_Saving_0/Interrupt_Generator_0/counter[5]_net_1\, Y
         => HIEFFPLA_NET_0_75248);
    
    HIEFFPLA_INST_0_55399 : XO1A
      port map(A => HIEFFPLA_NET_0_75529, B => 
        \Communications_0/UART_0/tx_clk_count_i_0[5]\, C => 
        HIEFFPLA_NET_0_75527, Y => HIEFFPLA_NET_0_75521);
    
    HIEFFPLA_INST_0_68053 : XOR2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        Y => HIEFFPLA_NET_0_72744);
    
    HIEFFPLA_INST_0_67868 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState_0[0]_net_1\, 
        B => HIEFFPLA_NET_0_72757, C => HIEFFPLA_NET_0_72776, Y
         => HIEFFPLA_NET_0_72783);
    
    HIEFFPLA_INST_0_67568 : AO1
      port map(A => HIEFFPLA_NET_0_72946, B => 
        HIEFFPLA_NET_0_72957, C => HIEFFPLA_NET_0_72824, Y => 
        HIEFFPLA_NET_0_72850);
    
    HIEFFPLA_INST_0_60944 : OR3A
      port map(A => HIEFFPLA_NET_0_74338, B => 
        HIEFFPLA_NET_0_74336, C => HIEFFPLA_NET_0_74297, Y => 
        HIEFFPLA_NET_0_74314);
    
    HIEFFPLA_INST_0_69197 : AOI1C
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[9]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[8]_net_1\, 
        C => HIEFFPLA_NET_0_72556, Y => HIEFFPLA_NET_0_72449);
    
    HIEFFPLA_INST_0_55158 : AND2B
      port map(A => HIEFFPLA_NET_0_75565, B => 
        HIEFFPLA_NET_0_75567, Y => HIEFFPLA_NET_0_75572);
    
    HIEFFPLA_INST_0_67609 : NAND3C
      port map(A => HIEFFPLA_NET_0_72838, B => 
        HIEFFPLA_NET_0_72828, C => HIEFFPLA_NET_0_72827, Y => 
        HIEFFPLA_NET_0_72843);
    
    \Data_Saving_0/Packet_Saver_0/state[0]\ : DFN0E1C1
      port map(D => HIEFFPLA_NET_0_74761, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => 
        General_Controller_0_en_data_saving, Q => 
        \Data_Saving_0/Packet_Saver_0/state[0]_net_1\);
    
    HIEFFPLA_INST_0_70439 : AX1C
      port map(A => \Timekeeper_0_microseconds[7]\, B => 
        HIEFFPLA_NET_0_72159, C => \Timekeeper_0_microseconds[8]\, 
        Y => HIEFFPLA_NET_0_72129);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_raw[18]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[2]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72280, Q => \Sensors_0_pressure_raw[18]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[1]\ : 
        DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72299, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72221, Q => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[1]_net_1\);
    
    HIEFFPLA_INST_0_69627 : NOR2A
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0/state[1]_net_1\, 
        B => HIEFFPLA_NET_0_72424, Y => HIEFFPLA_NET_0_72341);
    
    HIEFFPLA_INST_0_57950 : AOI1
      port map(A => \Sensors_0_acc_time[14]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_0[12]_net_1\, 
        C => HIEFFPLA_NET_0_74895, Y => HIEFFPLA_NET_0_74896);
    
    \Science_0/ADC_READ_0/chan2_data[3]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[9]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73419, Q => \Science_0_chan2_data[3]\);
    
    HIEFFPLA_INST_0_57326 : AO1
      port map(A => \Sensors_0_pressure_temp_raw[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[10]_net_1\, 
        C => HIEFFPLA_NET_0_74856, Y => HIEFFPLA_NET_0_75076);
    
    HIEFFPLA_INST_0_58322 : AO1
      port map(A => \Sensors_0_gyro_x[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_74801, Y => HIEFFPLA_NET_0_74802);
    
    HIEFFPLA_INST_0_58250 : AO1
      port map(A => \Sensors_0_gyro_time[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75112, Y => HIEFFPLA_NET_0_74820);
    
    \Science_0/ADC_READ_0/cnt[4]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73287, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73242, Q => 
        \Science_0/ADC_READ_0/cnt[4]_net_1\);
    
    \Communications_0/UART_1/tx_state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_75383, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_state[1]_net_1\);
    
    HIEFFPLA_INST_0_62567 : AO1A
      port map(A => HIEFFPLA_NET_0_73801, B => 
        HIEFFPLA_NET_0_73790, C => HIEFFPLA_NET_0_73954, Y => 
        HIEFFPLA_NET_0_73955);
    
    HIEFFPLA_INST_0_58027 : AND2
      port map(A => \Science_0_exp_packet_0[17]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        Y => HIEFFPLA_NET_0_74875);
    
    HIEFFPLA_INST_0_57713 : AO1B
      port map(A => \Sensors_0_acc_time[0]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74961, Y => HIEFFPLA_NET_0_74962);
    
    HIEFFPLA_INST_0_63486 : MX2
      port map(A => HIEFFPLA_NET_0_73683, B => 
        HIEFFPLA_NET_0_73675, S => HIEFFPLA_NET_0_73621, Y => 
        HIEFFPLA_NET_0_73758);
    
    HIEFFPLA_INST_0_62856 : NOR3B
      port map(A => HIEFFPLA_NET_0_73907, B => 
        HIEFFPLA_NET_0_73948, C => HIEFFPLA_NET_0_73810, Y => 
        HIEFFPLA_NET_0_73880);
    
    \General_Controller_0/sweep_table_step_id[3]\ : DFN1E0C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73926, Q => 
        \General_Controller_0/sweep_table_step_id[3]_net_1\);
    
    HIEFFPLA_INST_0_56913 : MX2
      port map(A => HIEFFPLA_NET_0_74987, B => 
        HIEFFPLA_NET_0_74915, S => 
        \Data_Saving_0/Packet_Saver_0/word_cnt_0[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75196);
    
    \Science_0/ADC_READ_0/chan7_data[4]\ : DFN1E0C1
      port map(D => \Science_0/ADC_READ_0/data_b[10]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73421, Q => \Science_0_chan7_data[4]\);
    
    HIEFFPLA_INST_0_66765 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[3]_net_1\, 
        B => ACCE_SCL_c, Y => HIEFFPLA_NET_0_73040);
    
    HIEFFPLA_INST_0_69916 : OA1C
      port map(A => HIEFFPLA_NET_0_72285, B => 
        HIEFFPLA_NET_0_72284, C => 
        \Sensors_0/Pressure_Sensor_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72267);
    
    HIEFFPLA_INST_0_61564 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[63]\, B => 
        \Timekeeper_0_milliseconds[23]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74183);
    
    \Science_0/ADC_READ_0/exp_packet_1[73]\ : DFN1E0
      port map(D => \Timekeeper_0_microseconds[17]\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[73]\);
    
    \Science_0/ADC_READ_0/chan1_data[8]\ : DFN1E1C1
      port map(D => \Science_0/ADC_READ_0/data_a[14]_net_1\, CLK
         => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73420, Q => \Science_0_chan1_data[8]\);
    
    \UC_CONSOLE_EN_pad/U0/U0\ : IOPAD_IN
      port map(PAD => UC_CONSOLE_EN, Y => 
        \UC_CONSOLE_EN_pad/U0/NET1\);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_6\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[10]\\\\\, CLK => 
        CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_6_Q\);
    
    HIEFFPLA_INST_0_56261 : AO18
      port map(A => HIEFFPLA_NET_0_75291, B => 
        HIEFFPLA_NET_0_75277, C => HIEFFPLA_NET_0_75341, Y => 
        HIEFFPLA_NET_0_75324);
    
    \Science_0/ADC_READ_0/cnt[0]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73292, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73242, Q => 
        \Science_0/ADC_READ_0/cnt[0]_net_1\);
    
    \Timekeeper_0/milliseconds[16]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72109, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[16]\);
    
    HIEFFPLA_INST_0_65633 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt4dn[4]_net_1\, B => 
        HIEFFPLA_NET_0_73329, C => 
        \Science_0/ADC_READ_0/cnt4dn[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73322);
    
    HIEFFPLA_INST_0_67193 : NOR3B
      port map(A => HIEFFPLA_NET_0_72957, B => 
        HIEFFPLA_NET_0_72959, C => HIEFFPLA_NET_0_72948, Y => 
        HIEFFPLA_NET_0_72942);
    
    \General_Controller_0/constant_bias_voltage_0[4]\ : DFN1E1C1
      port map(D => 
        \General_Controller_0/temp_first_byte[4]_net_1\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_74320, Q => 
        \General_Controller_0/constant_bias_voltage_0[4]_net_1\);
    
    \FMC_NOE_pad/U0/U1\ : IOIN_IB
      port map(YIN => \FMC_NOE_pad/U0/NET1\, Y => FMC_NOE_c);
    
    HIEFFPLA_INST_0_58062 : AO1
      port map(A => \Sensors_0_gyro_y[2]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75159, Y => HIEFFPLA_NET_0_74866);
    
    HIEFFPLA_INST_0_56288 : XNOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[7]\\\\\, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[6]\\\\\, C => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[5]\\\\\, Y => 
        HIEFFPLA_NET_0_75318);
    
    HIEFFPLA_INST_0_68175 : XOR2
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[0]_net_1\, 
        B => HIEFFPLA_NET_0_72714, Y => HIEFFPLA_NET_0_72715);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_WGRYSYNC[3]\\\\\ : 
        DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_20_Q\, 
        CLK => CLKINT_2_Y, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\WGRYSYNC[3]\\\\\);
    
    HIEFFPLA_INST_0_64948 : NOR2A
      port map(A => \I2C_PassThrough_0/state[1]_net_1\, B => 
        HIEFFPLA_NET_0_73518, Y => HIEFFPLA_NET_0_73507);
    
    HIEFFPLA_INST_0_69784 : AND2
      port map(A => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/ms_cnt[0]_net_1\, 
        B => 
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/state[4]_net_1\, 
        Y => HIEFFPLA_NET_0_72305);
    
    HIEFFPLA_INST_0_63365 : XA1
      port map(A => 
        \General_Controller_0/uc_rx_substate[3]_net_1\, B => 
        HIEFFPLA_NET_0_73535, C => HIEFFPLA_NET_0_73965, Y => 
        HIEFFPLA_NET_0_73771);
    
    HIEFFPLA_INST_0_60669 : MX2
      port map(A => HIEFFPLA_NET_0_74547, B => 
        HIEFFPLA_NET_0_74367, S => HIEFFPLA_NET_0_74341, Y => 
        HIEFFPLA_NET_0_74379);
    
    HIEFFPLA_INST_0_56453 : XOR3
      port map(A => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRYSYNC[3]\\\\\, B => 
        HIEFFPLA_NET_0_75321, C => HIEFFPLA_NET_0_75278, Y => 
        HIEFFPLA_NET_0_75279);
    
    \General_Controller_0/flight_state[4]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_74287, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \General_Controller_0/flight_state[4]_net_1\);
    
    HIEFFPLA_INST_0_62696 : NAND3C
      port map(A => HIEFFPLA_NET_0_73890, B => 
        HIEFFPLA_NET_0_73884, C => HIEFFPLA_NET_0_73781, Y => 
        HIEFFPLA_NET_0_73926);
    
    HIEFFPLA_INST_0_57933 : AO1
      port map(A => \Science_0_exp_packet_0[68]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[5]_net_1\, C
         => HIEFFPLA_NET_0_75129, Y => HIEFFPLA_NET_0_74901);
    
    \Data_Saving_0/Packet_Saver_0/data_out[30]\ : DFN0E0C1
      port map(D => HIEFFPLA_NET_0_75212, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_74763, Q => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[30]\);
    
    HIEFFPLA_INST_0_57494 : AO1
      port map(A => \ch3_data_net_0[7]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75029, Y => HIEFFPLA_NET_0_75030);
    
    HIEFFPLA_INST_0_67063 : AOI1C
      port map(A => \Sensors_0/Accelerometer_0/state_0[8]\, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[2]\, 
        C => HIEFFPLA_NET_0_72735, Y => HIEFFPLA_NET_0_72974);
    
    HIEFFPLA_INST_0_69087 : AND3B
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[12]_net_1\, 
        B => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[10]_net_1\, 
        C => HIEFFPLA_NET_0_72495, Y => HIEFFPLA_NET_0_72473);
    
    HIEFFPLA_INST_0_64367 : MX2
      port map(A => HIEFFPLA_NET_0_73713, B => 
        HIEFFPLA_NET_0_73705, S => HIEFFPLA_NET_0_73593, Y => 
        HIEFFPLA_NET_0_73633);
    
    \ACLK_pad/U0/U0\ : IOPAD_TRI
      port map(D => \ACLK_pad/U0/NET1\, E => \ACLK_pad/U0/NET2\, 
        PAD => ACLK);
    
    HIEFFPLA_INST_0_58070 : AO1
      port map(A => \Sensors_0_gyro_y[4]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[9]_net_1\, C
         => HIEFFPLA_NET_0_75157, Y => HIEFFPLA_NET_0_74864);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_x[15]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72553, Q => 
        \Sensors_0_gyro_x[15]\);
    
    HIEFFPLA_INST_0_69080 : OR2A
      port map(A => 
        \Sensors_0/Gyro_0/L3GD20H_Interface_0/subState[0]_net_1\, 
        B => HIEFFPLA_NET_0_72474, Y => HIEFFPLA_NET_0_72475);
    
    HIEFFPLA_INST_0_62216 : AND3
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => \General_Controller_0/uc_rx_state_0[1]_net_1\, C => 
        HIEFFPLA_NET_0_73860, Y => HIEFFPLA_NET_0_74027);
    
    HIEFFPLA_INST_0_66881 : AX1D
      port map(A => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[1]_net_1\, 
        B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[0]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/next_state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73012);
    
    HIEFFPLA_INST_0_62953 : AND3
      port map(A => HIEFFPLA_NET_0_73974, B => 
        HIEFFPLA_NET_0_73809, C => HIEFFPLA_NET_0_73921, Y => 
        HIEFFPLA_NET_0_73859);
    
    HIEFFPLA_INST_0_60832 : NAND2B
      port map(A => HIEFFPLA_NET_0_74548, B => 
        HIEFFPLA_NET_0_74349, Y => HIEFFPLA_NET_0_74350);
    
    HIEFFPLA_INST_0_58330 : AO1
      port map(A => \Sensors_0_acc_x[1]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[12]_net_1\, C
         => HIEFFPLA_NET_0_74799, Y => HIEFFPLA_NET_0_74800);
    
    \Science_0/ADC_READ_0/exp_packet_1[53]\ : DFN1E0
      port map(D => HIEFFPLA_NET_0_73271, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73243, Q => 
        \Science_0_exp_packet_0[53]\);
    
    \Communications_0/UART_1/tx_clk_count[8]\ : DFN1P1
      port map(D => HIEFFPLA_NET_0_75402, CLK => CLKINT_0_Y_0, 
        PRE => CLKINT_1_Y, Q => 
        \Communications_0/UART_1/tx_clk_count_i_0[8]\);
    
    HIEFFPLA_INST_0_55095 : AOI1
      port map(A => \Communications_0/UART_0/rx_state[0]_net_1\, 
        B => \Communications_0/UART_0/rx_clk_count[23]_net_1\, C
         => \Communications_0/UART_0/rx_state[1]_net_1\, Y => 
        HIEFFPLA_NET_0_75592);
    
    HIEFFPLA_INST_0_58190 : AO1
      port map(A => \Science_0_exp_packet_0[59]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_2[5]_net_1\, 
        C => HIEFFPLA_NET_0_75125, Y => HIEFFPLA_NET_0_74833);
    
    HIEFFPLA_INST_0_57049 : AOI1C
      port map(A => HIEFFPLA_NET_0_74888, B => 
        HIEFFPLA_NET_0_75033, C => 
        \Data_Saving_0/Packet_Saver_0/word_cnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_75176);
    
    HIEFFPLA_INST_0_55005 : XO1
      port map(A => \Communications_0/UART_0_recv[5]\, B => 
        \General_Controller_0_unit_id[5]\, C => 
        HIEFFPLA_NET_0_75614, Y => HIEFFPLA_NET_0_75618);
    
    HIEFFPLA_INST_0_66657 : OR3A
      port map(A => HIEFFPLA_NET_0_73132, B => 
        HIEFFPLA_NET_0_73071, C => HIEFFPLA_NET_0_73040, Y => 
        HIEFFPLA_NET_0_73072);
    
    \General_Controller_0/status_bits_1[44]\ : DFN1
      port map(D => HIEFFPLA_NET_0_74202, CLK => CLKINT_0_Y_0, Q
         => \Data_Hub_Packets_0_status_packet[44]\);
    
    HIEFFPLA_INST_0_65513 : AND2
      port map(A => HIEFFPLA_NET_0_73348, B => 
        \Science_0/ADC_READ_0/cnt3dn[3]_net_1\, Y => 
        HIEFFPLA_NET_0_73357);
    
    HIEFFPLA_INST_0_64484 : NOR3A
      port map(A => \General_Controller_0/uc_tx_state[14]_net_1\, 
        B => HIEFFPLA_NET_0_73559, C => 
        Communications_0_uc_tx_rdy, Y => HIEFFPLA_NET_0_73617);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_READ_RESET_P_0\ : DFN1C0
      port map(D => \Data_Saving_0/FPGA_Buffer_0/DFN1C0_2_Q\, CLK
         => CLKINT_2_Y, CLR => \AFLSDF_INV_37\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\);
    
    AFLSDF_INV_22 : INV
      port map(A => \Science_0/ADC_READ_0/chan[1]_net_1\, Y => 
        \AFLSDF_INV_22\);
    
    \General_Controller_0/sweep_table_read_value[3]\ : DFN1E1
      port map(D => HIEFFPLA_NET_0_74161, CLK => CLKINT_0_Y_0, E
         => HIEFFPLA_NET_0_73984, Q => 
        \General_Controller_0/sweep_table_read_value[3]_net_1\);
    
    HIEFFPLA_INST_0_67048 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0_i2c_addr[3]\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_write_done\, 
        C => HIEFFPLA_NET_0_72978, Y => HIEFFPLA_NET_0_72979);
    
    HIEFFPLA_INST_0_68494 : AO1B
      port map(A => HIEFFPLA_NET_0_72689, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/state[3]_net_1\, C => 
        HIEFFPLA_NET_0_72636, Y => HIEFFPLA_NET_0_72637);
    
    HIEFFPLA_INST_0_65711 : XA1
      port map(A => \Science_0/ADC_READ_0/cnt4up[3]_net_1\, B => 
        HIEFFPLA_NET_0_73307, C => HIEFFPLA_NET_0_73309, Y => 
        HIEFFPLA_NET_0_73302);
    
    \General_Controller_0/sweep_table_samples_per_step[7]\ : 
        DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[7]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_74012, Q => 
        \General_Controller_0/sweep_table_samples_per_step[7]_net_1\);
    
    HIEFFPLA_INST_0_66857 : NOR3A
      port map(A => HIEFFPLA_NET_0_73014, B => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[4]_net_1\, 
        C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/state[2]_net_1\, 
        Y => HIEFFPLA_NET_0_73020);
    
    HIEFFPLA_INST_0_67699 : NOR2A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[5]_net_1\, 
        B => \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[3]\, 
        Y => HIEFFPLA_NET_0_72821);
    
    \FMC_DA_pad[7]/U0/U1\ : IOTRI_OB_EB
      port map(D => \FMC_DA_c[7]\, E => \VCC\, DOUT => 
        \FMC_DA_pad[7]/U0/NET1\, EOUT => \FMC_DA_pad[7]/U0/NET2\);
    
    HIEFFPLA_INST_0_67854 : NOR3A
      port map(A => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[7]_net_1\, 
        B => HIEFFPLA_NET_0_72786, C => 
        \Sensors_0/Accelerometer_0/state[8]\, Y => 
        HIEFFPLA_NET_0_72787);
    
    HIEFFPLA_INST_0_56002 : NAND3
      port map(A => HIEFFPLA_NET_0_75371, B => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[7]\\\\\, C
         => \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[6]\\\\\, 
        Y => HIEFFPLA_NET_0_75372);
    
    HIEFFPLA_INST_0_66423 : NOR3A
      port map(A => HIEFFPLA_NET_0_73148, B => 
        HIEFFPLA_NET_0_73043, C => 
        \Sensors_0/Accelerometer_0/I2C_Master_0/bitcnt[1]_net_1\, 
        Y => HIEFFPLA_NET_0_73125);
    
    HIEFFPLA_INST_0_63806 : MX2
      port map(A => 
        \General_Controller_0/sweep_table_samples_per_step[5]_net_1\, 
        B => \General_Controller_0/sweep_table_points[5]_net_1\, 
        S => \General_Controller_0/uc_tx_state[0]_net_1\, Y => 
        HIEFFPLA_NET_0_73708);
    
    \Pressure_Signal_Debounce_0/state[1]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_73474, CLK => \m_time[7]\, CLR
         => CLKINT_1_Y, Q => 
        \Pressure_Signal_Debounce_0/state[1]_net_1\);
    
    HIEFFPLA_INST_0_70658 : XA1B
      port map(A => HIEFFPLA_NET_0_72024, B => 
        \Timing_0/s_count[5]_net_1\, C => HIEFFPLA_NET_0_72058, Y
         => HIEFFPLA_NET_0_72052);
    
    \General_Controller_0/status_bits_1[39]\ : DFN1E1
      port map(D => CU_SYNC_c, CLK => CLKINT_0_Y_0, E => 
        HIEFFPLA_NET_0_74266, Q => 
        \Data_Hub_Packets_0_status_packet[6]\);
    
    HIEFFPLA_INST_0_65224 : AND3
      port map(A => \Pressure_Signal_Debounce_0/ms_cnt[4]_net_1\, 
        B => \Pressure_Signal_Debounce_0/ms_cnt[5]_net_1\, C => 
        HIEFFPLA_NET_0_73441, Y => HIEFFPLA_NET_0_73442);
    
    HIEFFPLA_INST_0_65343 : NOR2A
      port map(A => HIEFFPLA_NET_0_73400, B => 
        HIEFFPLA_NET_0_73244, Y => HIEFFPLA_NET_0_73404);
    
    HIEFFPLA_INST_0_58682 : AND2A
      port map(A => HIEFFPLA_NET_0_74704, B => 
        HIEFFPLA_NET_0_74666, Y => HIEFFPLA_NET_0_74705);
    
    \General_Controller_0/sweep_table_write_value[5]\ : DFN1E1
      port map(D => 
        \General_Controller_0/temp_first_byte[5]_net_1\, CLK => 
        CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[5]_net_1\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/pressure_time[20]\ : 
        DFN1E0C1
      port map(D => \Timekeeper_0_microseconds[20]\, CLK => 
        CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72272, Q => \Sensors_0_pressure_time[20]\);
    
    HIEFFPLA_INST_0_61484 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[53]\, B => 
        \Timekeeper_0_milliseconds[13]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74193);
    
    HIEFFPLA_INST_0_62371 : AND2
      port map(A => HIEFFPLA_NET_0_74091, B => 
        HIEFFPLA_NET_0_73959, Y => HIEFFPLA_NET_0_73995);
    
    HIEFFPLA_INST_0_62051 : AND2B
      port map(A => HIEFFPLA_NET_0_73885, B => 
        HIEFFPLA_NET_0_73893, Y => HIEFFPLA_NET_0_74063);
    
    HIEFFPLA_INST_0_60819 : XA1B
      port map(A => \GS_Readout_0/subState[2]_net_1\, B => 
        HIEFFPLA_NET_0_74345, C => HIEFFPLA_NET_0_74350, Y => 
        HIEFFPLA_NET_0_74353);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[6]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[6]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72279, Q => 
        \Sensors_0_pressure_temp_raw[6]\);
    
    HIEFFPLA_INST_0_62749 : OR3B
      port map(A => HIEFFPLA_NET_0_73809, B => 
        HIEFFPLA_NET_0_73907, C => 
        \General_Controller_0/uc_rx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73914);
    
    HIEFFPLA_INST_0_64177 : NAND3C
      port map(A => HIEFFPLA_NET_0_73752, B => 
        \General_Controller_0/uc_tx_state[12]_net_1\, C => 
        \General_Controller_0/uc_tx_state[14]_net_1\, Y => 
        HIEFFPLA_NET_0_73656);
    
    HIEFFPLA_INST_0_57255 : AND2
      port map(A => \Data_Hub_Packets_0_status_packet[62]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select[8]_net_1\, Y
         => HIEFFPLA_NET_0_75108);
    
    HIEFFPLA_INST_0_70400 : AX1C
      port map(A => \Timekeeper_0_microseconds[11]\, B => 
        HIEFFPLA_NET_0_72152, C => 
        \Timekeeper_0_microseconds[12]\, Y => 
        HIEFFPLA_NET_0_72148);
    
    HIEFFPLA_INST_0_63902 : AND2
      port map(A => HIEFFPLA_NET_0_73662, B => 
        HIEFFPLA_NET_0_73594, Y => HIEFFPLA_NET_0_73692);
    
    \Sensors_0/Gyro_0/L3GD20H_Interface_0/gyro_z[1]\ : DFN1E1
      port map(D => \Sensors_0/Gyro_0/I2C_Master_0_data_out[1]\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72489, Q => 
        \Sensors_0_gyro_z[1]\);
    
    
        \Sensors_0/Pressure_Sensor_0/MS5611_01BA03_Interface_0/temp_raw[7]\ : 
        DFN1E1C1
      port map(D => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[7]\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72279, Q => 
        \Sensors_0_pressure_temp_raw[7]\);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/mag_x[2]\ : 
        DFN1E1
      port map(D => 
        \Sensors_0/Accelerometer_0/I2C_Master_0_data_out[2]\, CLK
         => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_72804, Q => 
        \Sensors_0_mag_x[2]\);
    
    \Sensors_0/Pressure_Sensor_0/I2C_Master_0/data_out[7]\ : 
        DFN0E1C1
      port map(D => PRESSURE_SDA_in, CLK => 
        ClockDivs_0_clk_800kHz, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_72395, Q => 
        \Sensors_0/Pressure_Sensor_0/I2C_Master_0_data_out[7]\);
    
    \Data_Saving_0/FPGA_Buffer_0/DFN1C0_1\ : DFN1C0
      port map(D => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\RGRY[9]\\\\\, CLK => 
        CLKINT_0_Y_0, CLR => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/DFN1C0_1_Q\);
    
    HIEFFPLA_INST_0_66249 : AND2
      port map(A => \Science_0/SET_LP_GAIN_0/state[5]_net_1\, B
         => \Science_0/ADC_READ_0_G3[1]\, Y => 
        HIEFFPLA_NET_0_73167);
    
    HIEFFPLA_INST_0_64565 : NOR3A
      port map(A => \General_Controller_0/uc_tx_state[14]_net_1\, 
        B => HIEFFPLA_NET_0_73552, C => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, Y => 
        HIEFFPLA_NET_0_73600);
    
    HIEFFPLA_INST_0_62868 : AO1
      port map(A => HIEFFPLA_NET_0_73778, B => 
        HIEFFPLA_NET_0_73957, C => HIEFFPLA_NET_0_73885, Y => 
        HIEFFPLA_NET_0_73878);
    
    HIEFFPLA_INST_0_69147 : NAND3C
      port map(A => HIEFFPLA_NET_0_72456, B => 
        HIEFFPLA_NET_0_72448, C => HIEFFPLA_NET_0_72444, Y => 
        HIEFFPLA_NET_0_72460);
    
    \General_Controller_0/sweep_table_sample_skip[11]\ : DFN1E1C1
      port map(D => \General_Controller_0/uc_rx_byte[3]_net_1\, 
        CLK => CLKINT_0_Y_0, CLR => CLKINT_1_Y, E => 
        HIEFFPLA_NET_0_73936, Q => 
        \General_Controller_0/sweep_table_sample_skip[11]_net_1\);
    
    HIEFFPLA_INST_0_57522 : AOI1
      port map(A => \Science_0_exp_packet_0[22]\, B => 
        \Data_Saving_0/Packet_Saver_0/packet_select_1[5]_net_1\, 
        C => HIEFFPLA_NET_0_75020, Y => HIEFFPLA_NET_0_75021);
    
    \Data_Saving_0/FPGA_Buffer_0/_RAM4K9_QXI[3]_\ : RAM4K9
      port map(ADDRA11 => AFLSDF_GND, ADDRA10 => AFLSDF_GND, 
        ADDRA9 => AFLSDF_GND, ADDRA8 => \GND\, ADDRA7 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[7]\\\\\, 
        ADDRA6 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[6]\\\\\, 
        ADDRA5 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[5]\\\\\, 
        ADDRA4 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[4]\\\\\, 
        ADDRA3 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[3]\\\\\, 
        ADDRA2 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[2]\\\\\, 
        ADDRA1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[1]\\\\\, 
        ADDRA0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_WADDR[0]\\\\\, 
        ADDRB11 => AFLSDF_GND, ADDRB10 => \GND\, ADDRB9 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\, 
        ADDRB8 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[8]\\\\\, 
        ADDRB7 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[7]\\\\\, 
        ADDRB6 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[6]\\\\\, 
        ADDRB5 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[5]\\\\\, 
        ADDRB4 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[4]\\\\\, 
        ADDRB3 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[3]\\\\\, 
        ADDRB2 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[2]\\\\\, 
        ADDRB1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[1]\\\\\, 
        ADDRB0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[0]\\\\\, 
        DINA8 => \GND\, DINA7 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[27]\, DINA6 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[26]\, DINA5 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[19]\, DINA4 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[18]\, DINA3 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[11]\, DINA2 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[10]\, DINA1 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[3]\, DINA0 => 
        \Data_Saving_0/Packet_Saver_0_data_out_0[2]\, DINB8 => 
        \GND\, DINB7 => \GND\, DINB6 => \GND\, DINB5 => \GND\, 
        DINB4 => \GND\, DINB3 => \GND\, DINB2 => \GND\, DINB1 => 
        \GND\, DINB0 => \GND\, WIDTHA0 => \VCC\, WIDTHA1 => \VCC\, 
        WIDTHB0 => \VCC\, WIDTHB1 => \GND\, PIPEA => \GND\, PIPEB
         => \GND\, WMODEA => \GND\, WMODEB => \GND\, BLKA => 
        \Data_Saving_0/FPGA_Buffer_0/MEMWENEG\, BLKB => 
        \AFLSDF_INV_1\, WENA => \GND\, WENB => \VCC\, CLKA => 
        CLKINT_0_Y_0, CLKB => CLKINT_2_Y, RESET => 
        \Data_Saving_0/FPGA_Buffer_0/WRITE_RESET_P_0\, DOUTA8 => 
        OPEN, DOUTA7 => OPEN, DOUTA6 => OPEN, DOUTA5 => OPEN, 
        DOUTA4 => OPEN, DOUTA3 => OPEN, DOUTA2 => OPEN, DOUTA1
         => OPEN, DOUTA0 => OPEN, DOUTB8 => OPEN, DOUTB7 => OPEN, 
        DOUTB6 => OPEN, DOUTB5 => OPEN, DOUTB4 => OPEN, DOUTB3
         => OPEN, DOUTB2 => OPEN, DOUTB1 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[3]\\\\\, DOUTB0 => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\QXI[2]\\\\\);
    
    HIEFFPLA_INST_0_66935 : NAND3C
      port map(A => HIEFFPLA_NET_0_73000, B => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/state[0]_net_1\, 
        C => HIEFFPLA_NET_0_72745, Y => HIEFFPLA_NET_0_73001);
    
    HIEFFPLA_INST_0_62609 : NOR3A
      port map(A => HIEFFPLA_NET_0_73905, B => 
        HIEFFPLA_NET_0_73890, C => HIEFFPLA_NET_0_73776, Y => 
        HIEFFPLA_NET_0_73946);
    
    \General_Controller_0/ext_rx_state[0]\ : DFN1C1
      port map(D => HIEFFPLA_NET_0_74301, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \General_Controller_0/ext_rx_state[0]_net_1\);
    
    HIEFFPLA_INST_0_64708 : OR2A
      port map(A => Communications_0_uc_tx_rdy, B => 
        HIEFFPLA_NET_0_73552, Y => HIEFFPLA_NET_0_73556);
    
    HIEFFPLA_INST_0_61532 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[59]\, B => 
        \Timekeeper_0_milliseconds[19]\, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74187);
    
    HIEFFPLA_INST_0_60855 : AX1
      port map(A => \GS_Readout_0/subState[2]_net_1\, B => 
        HIEFFPLA_NET_0_74387, C => 
        \GS_Readout_0/subState[3]_net_1\, Y => 
        HIEFFPLA_NET_0_74340);
    
    HIEFFPLA_INST_0_65886 : OA1C
      port map(A => HIEFFPLA_NET_0_73262, B => 
        \Science_0/ADC_READ_0_G1[1]\, C => HIEFFPLA_NET_0_73415, 
        Y => HIEFFPLA_NET_0_73264);
    
    \Timekeeper_0/milliseconds[14]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_72111, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_72091, Q => 
        \Timekeeper_0_milliseconds[14]\);
    
    \Data_Saving_0/FPGA_Buffer_0/\\\\DFN1C0_MEM_RADDR[9]\\\\\ : 
        DFN1C0
      port map(D => HIEFFPLA_NET_0_75258, CLK => CLKINT_2_Y, CLR
         => \Data_Saving_0/FPGA_Buffer_0/READ_RESET_P_0\, Q => 
        \Data_Saving_0/FPGA_Buffer_0/Z\\\\MEM_RADDR[9]\\\\\);
    
    AFLSDF_INV_33 : INV
      port map(A => Sensors_0_pressure_new_data, Y => 
        \AFLSDF_INV_33\);
    
    HIEFFPLA_INST_0_71163 : AND3A
      port map(A => HIEFFPLA_NET_0_71975, B => 
        HIEFFPLA_NET_0_75359, C => HIEFFPLA_NET_0_75353, Y => 
        HIEFFPLA_NET_0_75354);
    
    \Science_0/DAC_SET_0/vector[6]\ : DFN1E1C1
      port map(D => HIEFFPLA_NET_0_73190, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, E => HIEFFPLA_NET_0_73212, Q => 
        \Science_0/DAC_SET_0/vector[6]_net_1\);
    
    HIEFFPLA_INST_0_62140 : OA1A
      port map(A => \General_Controller_0/uc_rx_state_0[0]_net_1\, 
        B => HIEFFPLA_NET_0_73778, C => HIEFFPLA_NET_0_74040, Y
         => HIEFFPLA_NET_0_74044);
    
    
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]\ : 
        DFN1C1
      port map(D => HIEFFPLA_NET_0_72729, CLK => CLKINT_0_Y_0, 
        CLR => CLKINT_1_Y, Q => 
        \Sensors_0/Accelerometer_0/LSM303AGR_I2C_Interface_0/subState[1]_net_1\);
    
    HIEFFPLA_INST_0_68742 : NOR3A
      port map(A => HIEFFPLA_NET_0_72634, B => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[1]_net_1\, C => 
        \Sensors_0/Gyro_0/I2C_Master_0/bitcnt[0]_net_1\, Y => 
        HIEFFPLA_NET_0_72572);
    
    HIEFFPLA_INST_0_65684 : AND3
      port map(A => \Science_0/ADC_READ_0/cnt4dn[6]_net_1\, B => 
        HIEFFPLA_NET_0_73322, C => 
        \Science_0/ADC_READ_0/cnt4dn[5]_net_1\, Y => 
        HIEFFPLA_NET_0_73310);
    
    HIEFFPLA_INST_0_58584 : AND2
      port map(A => \Eject_Signal_Debounce_0/ms_cnt[2]_net_1\, B
         => HIEFFPLA_NET_0_74733, Y => HIEFFPLA_NET_0_74729);
    
    HIEFFPLA_INST_0_58539 : AND2B
      port map(A => HIEFFPLA_NET_0_74739, B => 
        HIEFFPLA_NET_0_74749, Y => HIEFFPLA_NET_0_74740);
    
    HIEFFPLA_INST_0_64698 : OR3A
      port map(A => 
        \General_Controller_0/uc_tx_substate[1]_net_1\, B => 
        HIEFFPLA_NET_0_73563, C => 
        \General_Controller_0/uc_tx_substate[2]_net_1\, Y => 
        HIEFFPLA_NET_0_73560);
    
    HIEFFPLA_INST_0_65982 : NAND3A
      port map(A => HIEFFPLA_NET_0_73319, B => 
        \Science_0/ADC_READ_0/cnt4up[4]_net_1\, C => 
        HIEFFPLA_NET_0_73276, Y => HIEFFPLA_NET_0_73247);
    
    \General_Controller_0/sweep_table_write_value[10]\ : DFN1E1
      port map(D => \General_Controller_0/uc_rx_byte[2]_net_1\, 
        CLK => CLKINT_0_Y_0, E => HIEFFPLA_NET_0_73814, Q => 
        \General_Controller_0/sweep_table_write_value[10]_net_1\);
    
    HIEFFPLA_INST_0_64707 : NAND2B
      port map(A => 
        \General_Controller_0/uc_tx_substate[3]_net_1\, B => 
        \General_Controller_0/uc_tx_substate[4]_net_1\, Y => 
        HIEFFPLA_NET_0_73557);
    
    HIEFFPLA_INST_0_61372 : MX2
      port map(A => \Data_Hub_Packets_0_status_packet[4]\, B => 
        General_Controller_0_en_sensors, S => 
        HIEFFPLA_NET_0_74266, Y => HIEFFPLA_NET_0_74207);
    
    GND_power_inst1 : GND
      port map( Y => GND_power_net1);

    VCC_power_inst1 : VCC
      port map( Y => VCC_power_net1);


end DEF_ARCH; 
